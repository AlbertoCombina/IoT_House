PK   �r�X8�uȇ	  V     cirkitFile.jsonŜK��8��J��Z^�Uԣ��,�9̤�,f�!KTZ;n�+��d��Ò���R���A��XUd��zM��V�n���m�e]yw�L����_����[�ռ��_�t��ݽ�o����~V?���V�1��0�(r�ca"?	���4
uZ(\����{x�����k�9�̑gnx�!�<��<�;&w�	�b����)&{�	�"����� 1��"d>&z᧡	}�q���.�\��4s�֬���k&��m��k&��I�fR���kf��̠����?`��t�����?`�L���0�C&�8�_qB?2�En��D��"]d��Lt������Ȓg�ܱ���k�f�c4�Yw{�?�ݬ^�s���t����E����bD��"^"/���D�:!xe�U2�*~��J�`%����dA�q�AC��F�b-C���2k���Z�b-C����Z&k�A�b���J	�A�b��d(�A�b��e(Ǝb��+O��(T�P�2��(C1�P�2�7)�9�]l��g�^
c������]�ik����n�&]2w�|/Z��xA/F�K(�%��xId��W�^%����W� �dV2+���J�b-C���2k���Z�b-C���X�P�e(�A�b*%d(�A�b��d(�A�b��e(F�Q�"��e(F�Q�b��e(6oR<z�����R���yq���~k�����7�&�K���|�L3����nr�xw��Y����4"���4�xq��q7�}����H�|hZ\'�s�H��z��"~�3Es�6����I��uQx�S�M�sϘ���%��f�����i2�#�}̴O������*.����R��v�?�ه{t�S�S��T�#%�S��Ts9�\N5�S͍��05�D��\����$�D��\�K"pI.��%�;�9����`"��䂉\0�&r�D.���� s��ʸjf�9�8�G�\�F?&��M�����_��p̘�C�t�TdQ��}�}�����o�	�t���HU��"eEڊ��+2Pd��Bw��B��&M�,4Yh��ddd]w�����������; $$$$$ӽ�:f�OG�n�$I��QE>�A�*_�:2 �*2�d�򉛕M?�mi.��+)p���e��]��zY�y<v�RX���a��ұ�2]�%M���y���M��`v"u)�[Q��P�\��M�E�6tW��e�n{^�K�7������_�K�M��M[Z� �LR�.����x@��Q��8qO11q�����Lc�1w}�<�E�;Γ<�1˵����s�� ɔ��%�����c�ԦU�u4&M��)���﮷Y��ɖv{����LL<N Ԯ�I���B�^���43q����1х ����v����F�I�1
jjBhsB׹x
H}�N�� 8����% =���&��O_ShH%�^h�Z8�>�`�n9V�
�w��s%ԺW���@^ �v�a5s�K��K��a����yݔE�%jX���0Q�k�Z&���F"}[w#Eɠ8��8,V�mq<��9Gmzq��̜�Uoʜ
 ��\�; 8�k���c���#ɰ�������hdP~4����V8��a�.��tO��&?�7(�8v1(	�"����*�3�n��n���
�#Ǡ$�8���瀹��� ��]����A��.��U���M^���婩�.9��R��"�C��x��p�Ec�.��@f\*���$y�.e@��*�*ⷳ訂�<�6嗧�"�:^)�j�<��A���p�g��{_??���4N{�6e��u�J���Nc�}M����_��zV��y����󻵭�u�6U�<y�o���l�����n�iS�ߏ�_�7ute�UN����S�:���t���M�bY������,ۧ�}۝���"����ԛ*�{�y۩Cg�u��K�}n�����*�N�|���־u�=����~���_��{]�U��������������7n4�~�/��w�����BW׹��*
��I=�D!.��B���Z��6?TE�֤+e�b�J��|�~k����P�f[�H�1��miMuݙGO	����L<ui��G?�.����U!i~;��~�%������/��m�����Oz�6w�3�{^d���v�t̼�̅��q����w����v�l���5n�ݹjҗϢ}s�)׽U]� ��O����l�ц�SqO��] ^�ջ�󴸞����0�
]�����Z��}.��r�g\j�9��㏙��QwJP�&�(A�AZ��X� �S�]�:�J�A6���v��i�pAj��o�I�J� %L*Q������t����)A�ZhF���Z?����S�[�ڦt5�K^�u��$�oi�I����]Q��u'�t�����Y�����\m���oPK   �r�X����7  �  /   images/2b66d102-ef9e-4dde-8ee7-817842500f7b.png�XwPS��� R���PBU�!��B	M@E)R tH�J�^�JGH�.ҋ�PD�@QJ	
�}��͛�����:{�{�:���={�8c]����dddtp=��YD��
p6z�d�>��zh226�s���v�^"������dTg	�E2�3v����3 �)������7?�s��ܒ�G��/�?�مg��EAFv�o�{�/�}yU��..��=��} �����ɋ	�F��>/��-+�>�1�Z�%��|�����p%��9�#|*xPݎC��S<�'���o�9�^>�W1L�Q3����.�Q��Օ_||�*~d �֋��'uy��j.��9Z�*� �u��+�>E�� �U�L�.5!>�n���f��f�q�7Q�>��-g�_�T,�X_k����>�:�c;����F+��g?���r�q�1�����Uʰ���r�S[0'H0]l��?�הۖrm��O�������98��W�8
�}�)��;C��r��3���&��?�.���d��ƛ�d��M��X�2U:B�72���/l�b��!�#8����G��d�{��x���m������#럀�(����ū�e��}��� }�g�
�B�!��R�����R��QD��z�_/�)��1@�2���X�L�d �IQ�l���Fb� ��yg�W�o��t�Cy =�(/O2I)IGP�yYr����?"yd�{n�y�kΊI���;���!����jx{����QB�
�����8/�<$���9_�B{���H��w���;�a���S����!EK��ű���"���l�4kf�Z����Y�5h[Y���z�_Q59:�eɔ��5
�Iu��qV}��Ԕ��� ����TH��.���F���b�	�mM@&�cA��	�)�����mگ��wD��M]�_����Z�)"�P��R3���Õ�m��~�y� ���,[=lo��� ��8,�Lć5��63�*(L|�H�	�A8h-����"Ҍ*{D��e`ß�Cy ��g\.�PK���$CX���U����a0|�.Ȣo����G��EE���Ϟ1�$��|�B�ܵ[֘hkת���(k
E=��/��-,�$bb�MLc�虅�/�6R=xW��4����ZЋ'R�Uf�8n$Ⲷ���5]P�I1ِݰ�C�d��{I��M�7��B�!�P%�A�ml�A��ƀ��$�R�zi�pT$5h��h�p�V+d��<�~`pn�Ȋ����	@7=*谭��x8-	�v�'4k�߲t�]�Eo��ʍ���\~5c�U��-�Y�Ԅ ���D���҇ӌT�L�%�I<�X�(�,v����Wn��L4����P69����'8�r�rI(�d���`�G0�G�14�k�:���
��$(�;���lEo�y�B��^z. Ul����i��n?	���L�{���S�1'�:����\ϴj����^P".�� �]�@�d����|�� [l�T;���|^^�+}T�{Y=мJ��x��]V=�IS��7D������o{_le�@x�0<<�e�R
@��Ʀ��I�Z��W4'Vc{Jq�Ukg��ʀ=?%e0W�-�TT=�	�!�fy{o�-+#*�S�OH�)� k�F�,ѽ3�L}k���n���G_�,}^]�Ԉ{|������yο-*7����U�j~�afh\��^"��h�!�`؟�l��?�g�MMc�|�S���X{7�E��!�����r�~��ۜa_�}�p��&��D��%q:��~Wh���05����v�7��Qskk�
Qf㦡!�og�%�Β��V��t� ^�kp���v73�E$��F-v^�.�*r��NbX�z���>r��y�5���+�9���9�֫Ƣ�z�x��]�@��E�]���z=�N����%~�.��"h)+�ѿ���k�7�W�u�����e�⹠�1�}�?��V�v�@g�Y�a������%���כZ���a{?pt�n�3�j2\>�e(oí��8�*��e��CU�sf&�����3�R�o�^=���ǡ�^1Q:V�n�z'B]�4"Z�\5�zH\ݭ�1�q\7�2�H�}������������O������a�	k��\�1������ȷ'<��S��VئҵJ���`��lu�f���tAK�a*d�$����f����V�8�zK֓�z�V_C��kj�g�^�l�A0e7��F�e(�͝�ga�5��i��ʘWk��zT0�MH�	p�۴�f�Fƭ�EFF�W�4�z7�P2[��`st�c��:S�@C$R|z��X��#OG^%�/)�vr��i�	>�v0ʓ}��S�U�+�Nf��V?���[�M�RG�;�]��m�mG������2��;��pk-ǳM>`���`'��X��wTtB���X�g�/�+�4��Ȓҋg�c�Yh���.��7Q�0?���U�S�zw9W��C%�6�u�mƵb�0�+Y����������
H�h2����*u���Y�>(iS�(�ɷ����4B��u�Z+��0�����t)� � ]�I�	KoL
�l�y����)���L�whm��<��-��>��=z�$��"[#b'��9!��r�������OO�h��u��vuᑑ~_��i�����D�~CNS�z�흟J؍�Pfa�~�ϊ�xUk�2�K�� K�U5�B5t�F��z�ќ�l�zO���w.�{�oj��1�xlb>3��b��F�4˸�i�D���k7��UT�X6=Dv�O�Z�2��LJ�94, n��P���L �}���mu�����d�o�K ��p�s+�`�z�gup��,ڒ�J����o�)��6��u��dw6��m
�gf?���o���<M7(p,�b7�碨��_��נ��{�)�d��2y��z�ɛ�-�2�1�g�72�"�r����k/��g���hA6�.*����T��IA{�P�4|>i���7=�%^��0d����J՞+����y�:j�I�h8w�OT�n���^�^N�s|\CZ�劻�Kp�zY�3Q�):��źC݁
��ƌ 42ji�*�}S�!�"����0V-ӧ;��e���:k����U�d�w��[\ȯ��dzzz�>���e������ Ґ#	�Z��N>�����R:C������@����ki�����e���j��1�F��\���?�J�<Q{�rO�����B�1^'m�����A�d�X)9qc��ai�w�j�gN�隄�>s
�\����24������5:��(Ǌ���d-�ޓ�=���rT�,@,d��FU��E!:S~���5|c^�-;-���:���X�)�4�M���*�0J4��n��Pa��o���\��g��ե+�z�[�)�o����Aw�f�KpK3���蘏�<���Fi���O����3�ҝp����,`-V��͊�5���EQ�n���y�!Rey)�ҵ���վ��9��j��*��v���j�Ǒ�����`���=�&��h����8��-b6m<�I��nq��9��Zb��B%��[��n^��l�%�W�۶��O�����)���pa����M\̞A_ix�쑋 џ���^�!��&''g!��x���">�V/���1�__��-H>���`l�;!}0\��Ee}ˋ�n�y��:f˻�j�)��� x5�K����u�pu�F*;p����%�@p���Hj�W�Q\����W=��������X�����Uݒ���J����G��ٮ��J��� ���DB�ʾ�����4ܡ/���%$s��5�N�fj�m��$�_RYu-�*3�gdd�J��l܋�fz��ʪ[��'d�U5;��td�_��?��ų��i4���� /5~��&b�.e�"r��R�2�Ƅ�A��FE]��%2δ����7+�,)�<��N���։]�ϯ3"�u�R��y�<����h���g��A�hr�ʡ�A�W9(�&D&��7���L�Z��$Ξ�o%C)�`0Sg��L��m�g��u�`W�ISc��W�|Lc4?!�4�ֶ�R��$U-=�N����g�r]�B��pq�ʒ�32d((0��B �{�,l%N���F��s�Cw����_G��^ʰW���ǜ������tsSl��͖�ҹ�q��W_=�[�	F<���N�5�Fc#�A:�J��ҩ�%HP_O_����X�����Ș�[&����y�n�-A��C����6���w�(y����N�a[�<i6��w(��q���Ige� l�4n���I���V�Phfӎ��8�tw*)�����Mӯ]y��Ap���*���#�������4��bq���snE��u	\�V�i�/PK   p�XE�U� z� /   images/3e05991d-8fe2-4671-87ec-9014655f7ce9.png�{w ���?)�a�"{Ʃ�CH��ʖ�%�8$['e���Ief���9���{�����wo���x��y����|<_��	��P�:�t����J��}r	�I�r�������Gw=HHL�Hib�IH���(��z�b���荔���V�܎0���k���5��M��w�H�C:�wde0D>���Ag&����ܗC�ߑ��G�)j+^lM�׎�׺��蹡t)).)N���bK������k���k!�n����Sڙ�_�|��f����}�g'�����Ӿ��0����7�0��Y�P�Ǉ���~l��5��G޺E���|��6�֚��=r����""с}I�����Қ�l�7���������ϸ�ͥ�y��̗�}j�;FN������=�׮$d&�M$�.�)��Q�S�(����q3�C e�)����}�g4��K�)��>����K�s�Ӎ/"�
q���kk���g�>��OǁL�X�O�,���ٓ����;�*Mz�Ro~χ�U�<�e�A��8����T��N�e�չ?� �@ƦwB��'�c�K�<��9�C���<�tvE�T���[�e�-@�Ib��ΡX�8L�H��$�}<�9}��O��N�p!sF}o�ɽ���X������ �`r�GP'��e�c�>"�"�_�P4q�˃(Ҹ��jK���U��5��1��wo��l�.'9|�7a���I&�Dޖ�$6��ɟ���$7a����*�z{9�}M��a�E�߭�� w�q3�����!h��$�����?�*p�A���^f���^�>~J�'�܈%�%���0)|)��ւ���x���B,��`c"�'y��[�Q�M�M_������ƴ'!렝��[��+���{(Ϡ�����*�J(Jg�Wu7��e)�`��+����i��O��`��}��|J(A��H�F3P�H"Ƽ ��V���������E��G@~��_}���]Q�JÛk�]ؓP�Y+�/{��c�����*$%�H@*����O'%q�#���ѠXݚ��\����C�W]^>�x7���p��&�X=}�����`>�}��w��O܁��u/��qs��l�V{�a�!��}]�i���}۞��}r@�P$��w�X)�t>��g�WV��Fu�G�2>�~��/4��_��DL������g� �*�V���RQ�
m\egZ �gJ��P�����S� t'#|��9\�y� �OK�K�B�c�a<�m�P�&�7Z�1z��⛁nv��Ys���a. qA�g�"��u 3��8��~��&���������< �2M�	�:�T�0��ҧܟDz������Ǥ3�Q��x�OH�y;Z9���)��h������>xB���մ�������pcǡ���h���,!_D�`w�k��.4��L���$]&�ʡ+��j�V���*��"z&���nn<���Qu���CTq%��Y���
A8�8+SD��$�3W�m� 3�@�t�+��0�}�FϏ-nMs;M�U/J���Q��`�]R�U,��P�1��AiLMŹ=�<�Q=c�]�ߜѷx?A��j#�46��A{�l������)ϫ�v�AԥM���V5�f���^�}�1��_�\M4o�R�8~�&����窈4��a���~�)��ؕT�Y�1�T��	KVg��n�!'���V��S�����p6��B��	?��W�wLi+6%�a
?����A�e~�Z� уh�>��
�s�,�XE5�4�I��nM��β�E������-.���'A�e�{�~{�N|C�����Mj]�#�#E�����
=nwd\�N	k�;�J
c��6�bOS��G��!����*�Ċ���2y�D8*.��m�$~T��<琅.��Ѭu/��*�$}�rA�w?b"B}�o����ٓ�%��LʎS�����,Ll�	*��t`�a �? x3�#��*_��=�{�y�a;���qY}��ۛ��=��@��R�;��L�� ��������r�C���d7��Z$}�!I�q����>.�T�5�?+p���G��>$AS��]i�����s<Jm�-O�m�P�t�&]3�����r<��O�TG���6��i˵Ӗ��[�W��W��"���; w��yF�狛��{��1�fJ�gfR�7��=5X�g
��fhz�w�w�ϒ�A�Ep���q�/�]�i��!�Mmd���
��U:�߫!ߜ�(�O�ĨN"�'3�L\P���M�r'\Z�-a���h����9��f|U�`�Q1�ɵ�&dw	�}�?��/11���F��^�D��`�z���9x��?�П_%e��������a����v+3?����o��{��� _����)��'o=��c�{JS�rp9(���=�]$G�?ؠ��!�p�,� ����0�?�q�QC�����2}�l&��Eoܑ���&�b�uO�����(e�as�E�j�T�8㣎Q�&?��8��^��]^�9zt%΍(��S�o��,.�~K>SM�5QjzF��,�Lh8�H�SQ���{-��ּ�c,ۣ{	n�Q�c�^H�ut���aty�;�l_
Ū����퐵�j��0�� w-	'�}�/�� kv���l���Fm%N�e�e ���k@��(�|]:�=E:�;��Q��_1�Cp������� ؏^N���sF��sA�߼#h.��c N�����Z�s����v���S^q�:J�%�7��GSsd����S^��
x�7��߸��qE��JY4�PG4��/Ɯ_���L=��哆����p[:����0K�9xR�2�?�A8�������b�@H��;��K+c�!�0kC�!�ؔ:o5��\{���"�D�w�5m�-��׼;,_/l��<`k8�<_�������+>�+� 3�m2����]V��J��$�ZTq����j��X�nnh�}:�'�ED��'B�L�@���!ErA�P��~���*f|��Ĵ�)�0"��`�UA���'�9��DA�R����=�KSoT#K�Ur�M�I�`}tu���-�KL17'��&�al�>����R ?�����d���?cfquNٍ�Aك�$�ڋ�z��0f@�X��<RW�G�*�F�c0�+��a�%Ŀ�p=�K4�&	"&�(�A����BRؑ8GZ2��_�wf���oq�/&���)�D��g� ��R�}_^�����V%���-�,6��$��p6�H��6-���u4���{ru��ǖ��7��w�	��\�
O=�z��pI�Q���:�Hʫ|Q���Ʀ<,4ZJl�9�����:S�k�j�K�9������#v�}���BK4.D��8N8���!�u�Tw�H��
���L/��=f�����!��1Q��AB
-P�$v�>��՗��[�m��A7Y���MK��N��]8�:/ly��e$:�C�ܱ[KIUn��?d-ʭ�}�,�/#�!>�c�uWXI�:ӽ��WV�F7N�Y�A���x�Gj�,f��M.�M=�e�ː��lFv�E�8� hq�9?U�=E����<aYǌ��00ܪ��n���$C&p6AϮs��a����I���Nq8�*R���e���	�,��T�"�+7� �)��c�����Y�B�\��H1���^��k�[]y�6]a9��?�X�b�fM���n�(��J�N,�����F�m/<�v���:xq'8�◘�q�~A��F/J٤����y�5����[\2[�%_G#p9�f�>���Hd��8؄=HrW�_��1��?�]��Yő�6�H�G���^*�A���=����6�y7����U�o8ywd���z�'ո!�+ke��E`ѠVX��3��5�����Ӎ\�q�˟O�����u�IWs�Phjt��`��C��IO��;Y6|dr{�*ϝ-�ʰa���j��5ڍ�[�5�lTZ\��*[����N~~-*��7v!�'ƹ���	����[�"�,юU8+O����bs��j+�Ϳ�k� o�s��B�Zo�)-��˹{��
e�ќȏ�y�9-���O�jz���~u\�)�/�/��:�m���T�ޣ8�O�N?\��nذm��2�M�]��;LA�۶p�ve��P��$�#
u��Uҹ��x������@%�x#B�T:�Dv���r�����F°(��⁫-B,���2��5��u�ۛ�M?�$B�P��e����+�~��6:��
�5�!�ʥs���o����l���;B:w"Tӳ�])��5��:�MZ�8
��5���j�p�ѓ��!��3L�	U��ݠ�dSb0ҶMJ�'��%B�|�zr| �x�����:��*���4�;�
���t��x��bh�9�r��TT~l.��F�{��y�A{K��pm�3�7X،w�>+z6N�W��F��Y�Vג��-��*o~TK��a���^kwB� 0��@x�x�z�Q��sLժ�{p�;���E�_���6%^�!Ș�E'��0}�H�S�0����g����(�	��oJl�8�lv}�D�����-���?�KW�) �����~�P�_E/��$X�6)��0��9iisC!K��̂�t�ŬB�	�|�q1Gf�5�ܜ���ڸ߾�Fjl�ad�,��< �.��o[��~I�p}��apV;�7��p��9۬'Ɉ�O��xT�v�t7�שc�c�&��~k�-�^X]��k�:u:��}�>�e�rԲ><�E�+��	7&Y����^���G�C~�ЎT����re�2� ��׏�PnL}�x�D&���͵�T1�,�����P�zC��6�W|>q���)S���3�4e]%6_��SN�en\�l�)�Kd��l*���z�D��5��������_�pV��Ij�W��d^�na8{��"Θ[E" M��Ev��\����R�_�������Aم�vѭ�=<]U�s\��?���\A��ߚ_K3���O{y����v�L����Qп��x��E�R���u>�6U����5ί'N�.��}�#��%A��J[=Ϻ5�.���z���\A�K�_�3���@�,M��Ɖ���O Z��|X�{�M |����KFcL�P�eF2��b*���c�_(3�B����4kNe�_����ͽo���Ku:O̕���5�G�E[GS����P��!J-��5�V�k�������i�J���l�����$�a��B�n� Q���[m��a���t	�F��	�~{Q��^��|I�0��(@|o�WՊ0���0MfI�J��v^����q62�Ԝ	@�$2��|��~�:C��_	7Ev:��\ö�H+[����D���cYu�{><��pS�݉Ӽ��1ϝt��,��9��&ˏGu�	V�y�,��48�W�8�K\��WL����,��4�9�3��D��r��U�G!�-J;:�ӼIɔ����v�T}YU7�.��~������ ?�+c5�M7i��G����Q���˚�w��v�R1@����`p�O��0��v�5��)<���_��t��sf���;V������@�DH%�j�jLh�j?�4�&	q��E\d'�.�}
�/[���VL���k`��։�P��y��&Ll5�����Ɠ%��
�-wY�?:FN������Z*��뻁��<��g��:g��1X ��4w�>��.��۟�<n��v��#"�6`����1�B^t���s%Åz������f�|����X�¶`��<c�X����c�-Ya8�gY�b��M	��w�3z�f�sN������~f���	���x�'�e�2�l���ދ+��
���(R&B�~,�pfi��E
��	!�$���^2B��5:��r�U�͉���a��ng�=Vݫ���c#�ݸ|��L��D>�?�uH��Y���:[z��Z��wy ͊��ڋ��;�*���M
'��a< hʽ�u���H�Sx�]��w��&�h�F��@
h�w�~���fJ)��Om�>Y��.Ĝ@�S�nx����(����J����c�ڭSS�d�.LJ�dd��u�gP4*!��*�:ي�� E�Ge}"h��� >�--P����}�E�G�i�ȶ�����z��*]*�;D���NѸ7���p/�Q���8��WR)I��>k�}���>�	D���R�f��Јo��%�����)�@). �*kP��Ԋ��3�V�I�W}��>\����v�I��N#]-�s�4b,��8K$B7���{de��
[E�j�["��</s)�w����=w��=V-�ue�HO��MW93������aH�]�u�B"D�:�uibj�Y����jNfw�G�=����X�K����d�|�� X�s=�X�K�}�`�v8�μ[8�v��c�#�(��N��1��Ŀ�R{dCE`�<�0v)�C�{W8���qoѾp�%A�PW�*W�x7i��䉒NI��k�Br�[��� )v����y�<k���Mk���-IF��[/�G��]q���M�P��o����w��i������
�W�6���or���� �i�j���`�����ٷ�bÊ�'X�ѧ�+H����M�y#
�zfXA��'���D��� �vbǲ��1w"X�k���-�\w���w��B�Mk."���Ң�}�D�]DSV��؄��$'�P1�Vy��i�,׸�~�FWe�h��$�߂M]o�uk�ٹ�S#��|P �8�4��o~ u���vt��ޓ�0���$�פ@*l��`�AšB=5&l(zRGW�訄`dd`�Dey�:�{J�q�����eL.t����A}��_��t07Gmh�FAGg,�F�������"� 8Ϟ����Q�38�w��0�}@�^��P�����r5�G�|wǷ����:�����7z�R�<lY7�3�hت�����!6�T��ݗ�bǿ�R���53����-��E�b�޷�2nUKݯ`��!�%��<��?��d��A�2�w �e�x<g�""'!����A�<^�x�Ŷ��2-}��z=S�W��C��D��qm��h}A6c�6���^��H�ڛi�MʈN�D�St��{�3�\(�0^Z����Ů��X�U��"��ܼ��P����-�}d;�fʎ�^�ي����h^��u��)!�C��Nqz4Db������)�
h�-��U�/��q,����N�^v�<�?����P��\���K�F��K{0��bW����]7���a�o�C7�ߖ��e͋z@��œ����;���s>��-�sW;$l<�@l��u�l�MS �p������A<��,YG�jb?��:ĎA��U��������<�#�bi�|Gۢ1F& ]!����C���5��ڙ����7�z�� t�=f�h1�m�z��ބ�3���n�ڛ���F��^�ղ[�"Rۨ&?��i�]K&�z̮��i۫n3�ǌ�e���ul�F1�VBVW��lS }�Z��W��{ ��9��ƅ�t��(Mt��*]ewr������]S|ĝ�.�= ƨ���Bl̐d&	G���殜��F׮Q�4r���N�bE�"`~s�G�_%�3C�=i?����g$��k����o����]�(G\\8V9�\��_��ŉ�7�Z�"�m��&�W-�ι|�0�5q� 3,�i@<�I���x�öW����AH�͓'`�|
4�^��Q��ts��"�q�w����:˵\�b�d�x�`6=�Q���ǌ�a�%�sא$b��Q ?�m��1���Uf-���S�x`��q�cdA9�id�L�b�v�h��l,GUZ��ܼ,�(�����l���iI�Ԍ��p���E4�����d��t���6'�4n�� #�G�e)T}�������D�ݛ���Z��q�Ql�yݲ��V�)kp���Sx�=G�{�୸�3�N�������3�h�s��~PJ̧:As���;�UN�S�������?�,g�]�G���82]�Ǐx�\1c �z�˘�7���ސ���#�����b<�,���Ȗ����J���X�x~��&��&��6��-�`հ�P����Q���Z��Mkl�"E|y��c�t+q���؇E�I�t�|����-.��	#JA��nɔ;|�{��ڷ@E'JQ�U#L,�S���Z�_�d"����Jqd�2�Ӛ�DS���%ٯ�\��Ѿ�p�@���I*uu�=�[>�"��蔇���a��3����ߩ_��웞Y��a6-����1t�t�Run��}w�/֚��:L��."���z'U�g��0��"ݖ��k���#��1o�Þ�~���O3���:FH!�m��X�K�uތ٦f\\���]�VO[�EÏ��#Jb��~lO�]��>-C��}��ې�>����S� �Ϋ���q�ěC��/���Z��:���:�I�=w�x<����-�j�>��={"���0�x�����C����e�=c P^��@v�����8ȝD��$��ߑ���Y����M�5����t�+�Ӿ}���k�7m<sX]�2� ������wA�:Ouʖ��R�Q)qG�ƛ��Y;J�������a��\����GНw�%`��ƛ�� ln�/�LLR<��l������)���ӑ�%�RM]���.C���Se$\[�q*��Л�%4�?����y�$@�x���	�āV�8m���D\�����|���ؒ���?���7. [<5�D������.ʐ�U��Z�$+S�]��rŞ�!�}��z�/��&+ia�U��]5�8�j!Fg�:F�f ��5�M#�xW�3�]h��*!�OO�I\)��ת�)�i��þ_xn�BJ�������-P�˵�cQ����Ҟ��[.��
I��vw�Cɨ��S&���$��j�Pt�+����@+[;�T'�����Z����%;���#��O~Β�]/�����;�����ß�+5��O��7������92��+ȹS��B�4	9M"�x\�l{0#0K�!��2�U#����A�)��;��Њ
�W�������ʛ�6�k�`g'���-�φ�?e���u2���=�����4Y %��Nn�Eh�.��wHQ�&��\7��nu3z�xFSٸ)鲊�X἗s��?�Q�~E��
�9��IK?fː&E������#�������@�Q�^�H��+� �",����t��4+�\� ��Kp�]�;ؑ��>tkg������o�43j�u�1(ޓ�S��G������$�֡�|�4��$i �Mw��t�TRkf���]��-}�?U����
�g�o�w��~��������	s���G<�6ޭ�q~���+�E	�g���u���[��cxg��U= ��W�}is�))=kI���8��#�᳨9m<x�'Sr�6��D�M�#!��%��q��w�k�Gv|�~|���4-���"0&/g᭭Pf���׎�}y�Bs���T�*tup��T�,�=��~./ ���QJ���2-V��)S^�˕�'��_���x�ߣ��dw�?�R����R���3^T�ԩS�H�����}�?�gAe�@��C�/���/h<�s�+`Z�
�[~��3j�TY�=�e��F�� � ������MJ�;���Z�*��a��Ћ��mL:�z.�j��ݛDg���	���q��Y��0f�[�l[��<�"W�1����⿓��.|�����xL�[n�h��qc�_��	M9�e�z�W��F�V����]��tC�)�؏'g�,�w���)��*d�����n�s@��d�"/�p��w!k�	�,�l)j9{r���Ծ��*U�46��$��	�n�}2�B����� ������ĤӈXJ0	��-{N�w5��d�>�HE,����fLl�X�@���زa�ɗ�q�R��:�����A����#J����uj`/l��A~G�y�C���0��a�n�.���|��P�v��R%ؠ�L��7�u.W����Hb_ƚ��&�8ɆW��=|��RB(/1�0U�ޘJXLʎ;.�m�?����g"�J�ؠR����bs����ݾ�v�S�]+I5M��ő��� mG���v]�[�I��!����1x����6��VT�������$޷�����p�Nn�O#doE>5���S2���z�]h�����H���KtÐ��ty^�֌��K����}�� $��I���z���6��a�Ђ�Z�a��Ρp�9H�d�u ]�����>�OO!b�M��6'v],ǂ�o;8�u��O�*:,t��0���,�b5B@8�5�\{�:;Rl��m������y�o+�{���gg_�y!�m��Y�U��Ҟ�_���|x��1½�s���]V��2D���ևE��r#	�����-����m/��������+n�kꅎ7�'�ؙC?�p�&���nJ�Μ�7+��`q�^�9��/_s�Zc��^��iјz���H��	�w����Ȫ�΀X�@WZP5���j��e{�C��*9-N�te}���l��$��6}3�j�ߴj%p��|8b�7p�c����~]8!�m��Q��.��J�[7�7�*!��j���;dw8������W)˞��C��K�M/��z@�����)��^/�=�e��ռ,&E����a~T9��\�I��R�L�ь>�<j�N2/���N���/@�k��:�9����v�z�*�6�`iز�����\�p:��SQ���?v��������JvE�%�N�ۮ�6�G�j</E��Q���l**��j^:�0͍J��:d���Lu���ES	e��(�3˹]��8����r�Dɩ#��ݛ��^5R��>:"�ˋ���u� }��G���;���}d�J+�ӎ^\L]n���w��ݻS}����io ]"@%&ړ��ഷ��'�uZ�d��|��;z"__9XX�[�M��0>��0‏��kɻm�mb�z�N?��L5�er������ڭ��d{��+~bw:���`�A�5IL�j�a��M;�����i)�i�HU�~���VW^X\Z`w}�UVY�H�����3���S
�����w4�Q����#xcs�&u-_s��_�ۻ�8�~��2��[a�Ud^��`~ܐVe�p��G-�j��6�f�a#v�k�7e:Fxi4\Ӏmk+Z��6W��|���"���w.�A�'��4ŒȘ�]����AZȂ���K�,Gu
.>n�����GB�5i�T��	�����Zs��vs���AK��B�>!
��>r=��a/�b?c2��}n�eU������T����yc�z	{��ҭw��MK���s��B��c���R����H]Zս�;��¾�{h�<�O7�� +.x������m����Rr2ǝ̣G|��qv:қ�#�-��L����T�͊a�����辩��ˬjy�'��MW�O`�d�_u���Tސ9�:���Wtآ�p﹧��0D�im���S����	��K:L�)C��m��z������-ҩ�R�R�][u����J�K�H�~���J��ÌF��]�|]=_}gɐ,��2���K��ĉZ8X�"�HK�p{J0�Xw�9�ǣ����0�V��G;���t�����U�o��!9�����O�^�`�nsk<֨\���z��qĻ㾙�}`���q��Q�ѯ�q��Fo�W��Mq��ꥌ�ź�l��~������ns��*�� ��wJ͈cV�*S���"=�����D�ٜ�(|��%r����<D��%�G�&����8������K/x���_P�~x/=���@��G�a�����G��jʫ����~þz笚Kܬ��o�Kޔ�u�y�6�ͣ��6L�6M�q(U���\�&��k�A�n| ?@HM��2�= N]��#��7�Ĝ�E�)8�}k���O�q8����v��H��^<;���4:=�<�lf����Eo-��ý�X[h�'��G�W�Ȃu/f��
WL��>�VB�ӕ�^���/q��Q5�����2�W}�Vw0�Liqmz�h�j(:�x��%�M:5�[X_�
��ъ�Tz�FvX�k��>]����#Kj��)h�����$o>�����'���뎚%��l���&Ǜ}]'�r<�/�\���A���gk_�pRɡ"�ƻ~�I�6�4���x Q�4��J�hؔ� ��1�_�u?�a
��a�R�d�weۻ_߈�]��e�;�m`��V����^t�x�|6z�����:U��лh�չo0]�n�.4�w��ڜ���[�A��U����<���PU�6���vnN���)y��j"K�-ix���.*0U�t�M����Խp�f�NA��`�ϔcS�L�k���v��O��=U���K����$��-͜k�3�(��Y���[�/P�<$镠m�d����yRP��_qNQ���k6��x@6{A�"�Q���8GJۇ����L�b������Y����v_�_@<а����vu�z��Q���E}l�n��l����B��81u��V�m���9�Tzi_ǢJ�pT�}zf�`���螐�KF��JW�'�p�'Y��ۣ<��N�v�:��"�c���������Rj<M ��e��Wn)�f_$!2d�3V'�<���㚶�����h*3��ߖ�nO�ᶠ�s𫉐51��T�l
��q���b�m�ن7�ä�gM��U��X�ZUԂQ/�hz�\w�|Ui�7t����r�F�q��6��w���O~������>_�6[־���t��^������(��
R�o-|�[��@J�A6��HV���t��ٻͻq�e���q��(�Q��$�Ю^$uo*�V�6ŏ�]��'2I5�*fJ��W�g>T��z�GY}=OC������/q��ۗf\�ϤI1���߷�.�C�4O��}a�~H� h
��a�&����	���C������Yʸǖ�?�0V���`Ii�R@��-��o���Uf�TўYǝ�*��E����)���zDr�]~!\<�v��s���O<Yp����afW�*3d�fM��5VI�Nf�H:�e��U�J���舉� #��f�NvX��U>�U3zU�BF�iՇZǗ��(��e�Z�>}|��-�o䪽���*��z*�� l��g�8����;�Q�)�U�lTM'iߧ;ҷ��U��5��w]*CD�u)|
B�j-k��1,�n��T��Xp=y|M}����3;��|��P+X\I�[5�B�hRm@���͙�ugr�-a)���Rh3�9t��Y	�`�M	�6�ȵt�'|��J/�K��Z�!t��;�Ǽ@�ȕEM=vϻ���v�X'��ǲ�{�4�@9��KD<EEF�G��N䷗6��o�1���K��5܋�`���JG<6;�q(�:1C���/��5�a�Ó+�i��wYA�%c�no��f���X���+l_X��KK/I&��u�U��q����p�|4��4�.�昉F�`�=��
���2����\86��|�G6�Jj��vl��4i�p�n��W ���s&B�س�����G}l��n�O�3f^+��A�R`g�`���u(y�!*]Vж���):�AR5����E(�Jò4��#�n���Ne�����DL��d7�w\�<���ᠦ�מ=�n�J}�A��w�ѠB�8�ɣGf���q �/E�v�n�A{ͫu�PʠX�����c�B��@�� V��AVun�Ѩ�����J+ߎt��!,�p����(������<�Y���x�L&�Ny�]irٛ0��U�e��6�I�~�-�ϢU[��}�7���N�����	y��p�*�a抉:�;�4J]�@�m�E1�#��o���-���~o4��,�$^�.�� yǁX|���Z��J��3��]{���&��U�n����L��A�C��/�r����+�d"e @���>e�8���E3�� �F�[��y_ׁ!�R�n�w3�����ݾ�va�k���M�;�h��s�%�]x�OE�#2�?]q�I�OT:P��fc�zk=¹
ϼ;�|�����]�7\>�
�X��/�h�C"��A���8W�hVP��'�U������ߗ�9��7..��#�g��,=��v��B�_옑x��9Q��;|`Ag<Ȳ{��]�����������Uμ/Y�;d����Y�/Ç��[��t'?)�F�.����,�=A���vQ�(w���mY<��-��U�T����g9�K��gEe�.�n}'���}��@Uٳ��Joߐ�Ϯ`34���k����Z(���h9ߏ�7j5X��.����d�}h$�i5��U.���W�TWrC���Yc�	K�X��̈́ơۑi��^9��j�����єݕ���`t\Ѽ�����G���ap����^BJ�&�.�u�y��0�3���]dz%J^�����r�R�"J���ZmN�]5:�ʃ�,����[�{����l \tDm��U�m*J�l��XȎ�&0����w�����|f!��T�v�ڶ���J�Uƽ�g���� E����nx�M�pm����SvVQu~Pf2��8��4����=G���}��j�����z_e��L��%Л%0��Q�Fu�o?�S�N�^Xe��+u�B�P��������Nz=�N��)8�q�wO�H?��u'����Ņ�=������'�l�ᦃ���֬�

�ɇ��B����ڣ"��#^֟ڱ[Q�|��u�����roH�F��?�L�>� Q����!��1<��}����`Z��N�x�G�����U�mM!�;v�ݜ'ZdC� �i~-����M��.=S���e �n>���ǿ{��Bud`��B�B\��:�l���cu�ϔ.78�P�˅d��5��ie�[aZē	����}TlF�;٨�5F�'.,��ڃ��8~;�GUkdkSg\KF�u��	�����t�(0VmŎ�Ixz���g)�Y�{k��N��S$/�J-�����M��������v_�^r����a���b~nB Q�k���	8Ry���m�_��V(85AmPr��5#�]��'�;��*x��%A��`w��7�C7+�~$d�ËF�72<����50�1c�Ϻwp=Q�9��ϧOb��F�G5Q�=y� �_q�26�m9�4��������.� �qYj�E�G~�/t��\oi�_ԄU���mo?���x�!a��A`��ň>�P�b�~A�*#װ�Cn��J��z��ʏjqs�R�!��� ���H�xb����>�3#:���<�4aB;�t�_�H '�8X�60v������hl�Fć4_C�te�ޯ3(��	m�M��L:�q�ۙ�(y^�t�� z��2@��@�I'��6Sz����yP���U�-��^���Q�򣞫�Ё�?�l1��3�:����<���V��D���b�ؿML�zI���;d�g�wlr}��|_�׉�{¹���W̠���'�ss��F*��̈́��U���[���Ef�RW�_D��쫟F��S��~)���=�$V����붧��M�zf����PŅe1�"�Z9k����&hadu�Dt��]Q�Y�=�[<��m��I��z�۞<��)��e��o�R���iMTN�@��@�jPj�S��r�Y��F�����ee���o�7�-a��,�T�߉~�d¡he���"���Z�bp����%�	G=>�h.�L^yE�-q Q�"]~����]���v%P%�չ�r��0�Ljqu�)��+�W�9d���ED��QuqKt
X��c�K�#A����|�0V�z����k���B��W��&-�{_9«������ě���Y��c���8��O�
��g���\�$��.>�y��j�z��I[H/J =���a��)*���k�1cU��V뵖ڃ���Oқ���K1@�7���Vøx�k����߇.�cد`;ۧn%r���������䍽�a�G����'��a����&̂Qa�8{�VH�h~lL�~�Ž�S�2p4e|��1�&T8/�5-[wS�p�G�i)��֘H*ȱvm�Zp�E��͹�qz�����e�+t�YJ�����խs���#
tZ'�+ZCN	G��6p�{�f��wZ$�M�����A�V����_g@�ڢHԿ���z4��,�u�_��Ŭ-)�u����!�0�{�4{K���Q��Q�Y���h-�V弦�+a�LLD�����R`qIz?��/�Gi��НCL������فk䁌����V>,�;��*(��"�~����|��~LuY՞r�8�ve�\�tQȐe����6�P_�S�1�kܓv�T���͝5Q�s�d!E`W-�A�YQ�=���L]�Տ�w}�����&�Ѣ��4+��!���S/�h��s֏^���a�H�/�Ou:QsK$�3����E�7Y�N���8����ו�45��	�R�-Ԍ����,�!�M� �e_� 3����o��pY�оY�O��@���)2����P�-���S|a�H�b\�8F������e��3�SS�ò��K�ϧEit�8~�ys�q(��8��r_|.Ǘ�*F�۝������l�f�ӕ�fL;3��������	n��E����RZ����d%��4����3C��'o��n����K���uM��f��s	���zӾ�Q�Ekn�1�ؼ��.���za��~p\�C���:�}�4�;��!QH-�t�Ad��,�F�_8Z4�螻���1t��]So��e��r��;�1�p,chȾb�X)˔���S�������#�f!����v�q����ӷ;���Y� N���gԼ����.͸��x֫I�]v����^B�����t��lg��~O1�8R��Ȼ̆D���.w�wp/�\ӠIZ|�v�����y2����(q��r�����R2r��Og���[��?&n�������� %s�:u�9k�Zi�+��-�:ҟ�0��4��F<d�
7C|��ߪ�����/�'/�����ߌ�B�*0����;\��6g��Q�X�]��0�0������Y�����O�@�c|�G�v@�t{��㲦�G�+����.����4�$%<�{J֧T���J������q�dک���2&P���$�L���.Wz��݉4�͢��}w<���!렒}i��G"E���W�8q��-dg����,㐽��9�98��>�;��y=���G��u]��{|����Cy�G�AYC��� $�x,q#�8v����E!�t�.AK�N*�/)pz��X�[��{6_�p�M�
$��p�n���ҹ�J�?�>P>U'�-�0�z�;M{�W+(Qc*d�-�@������r~E��*�b��a�� g�O"N~Nn�U����<K�*ፄ##
O�Λ��_�Y%N��]���v�Y�EIM�s�ƺ�����B�xb!��k�K��"�g��c��c,
��<�M��&��{�jK�*���ֹ�=��t���֐^�c:��NZr�����!O���K��OY���������˳�>��U�j����'��s[2�ǾV�gm�MӢ��4N�%�\��tCt�X�PQS���i����h6B�b�c�]�1WY���1�j��Јb�7<ϕ.�	�Ppi�C��of�XW��%�h�h��η���7�qX�����Q*��<�/���v9D�-��	n���r	��=�A��>@�7���ڮ��gR��`�1�S�o�T���*x�$��a�����vHQVK>-qHF�u�4�W�&��BЪ�b�l�S�A5?���qZ���>�զ��\>*t��g����AnH`Tǿ�P��gn�ypr�������F:�N��UO�*)D�����l7����Wy􊯻׈�7b�J�VƯ��vA�6��(]����uU���僷\2��G��:�����r�_tn)A��s�X�d�C}��9i�)��)�K�"��ߕ�x��D�La[�=��P��.�yƇ��-��HZ����zپPNd�ˌW|\�V�<w�����r���B���D)�,��*?���\XL?[��u�{��f��a����$���3;mq�A����֝|��EM#ޘCY��5�-��x2_>r�^�t���x!�8q	<�N�݄�+�틬��݆�fo����/H��%/�_��=�ꓸ���k�tmX�oS荣��[d�����kZ9F��J���D��|�r�C�`�ojeS�"Ĺ��/V�UK�)Z��͑�]�sDN5����N��Ɗa��p�����aY�FRzl�ל����ۃ^z^yF��3t�FRvM�$U��<	��DX;->�d��_g�e8ݷ�7��eCEK��u��递|6�i5�h���0�=�H`_�	B��y)VY!��:�wA��ɧ��Ns'�Ā��}&���b̾����/n}
��5���JZv˓EDH�J$�ړ����x�yl�x����;�,y⪩���a��/�m�c7]I�y�|��m��7�v���ɫ>v�뙙r`	e�_�]	e����X{�EL��#3�#�#5������s�v����ۏ���gWi[[�����X�5:
�7�x��=�my|E	�X�U��2w�g޽:Bo\�E�ۏ]�r���s|�x��b�����V���;a6�~��.`@��u�����W����6YY�rBg����K��Δ_I+�,x�U^�����=�v�N����5��b�����I���:�a��P��_n*���ؔr����{c��	�h[_���^�+��t��g���~�Q�_0��VZ}/���'�Ѿ|�xu��A�k�Ys��%�LQ5�f;W e ����|�
V�%
ZM�:��砶��|\�I�	!�&k���t�..����\�+.qz�k�Q�HX��[���C��<'��hp< Lc���-�K+<�ud~���vf{D=6F��ú���>t�%oG��<>����v�	̸+����L3�B���
 ��
��ٯMm�И�M��.�axI��v��:_�6��k�r����IevQp������j�[�}.i���E�U!�q^g�ɯ�^�|eHK�AbD)Wv�U��~�aX��v��ĻBi�˻�Ƿ�6sT����l��ި�$�G�p4b�/��)��mZU��Mζ�Υ���xf��(Ú�����Z��>�	��T|j��i�d��B�����T�%�/�������?����1Ն�;ü�#5N$G[@)f���������9��&[>n��`�'&Z�t$Z)�ߔ�C&�u< N��;��P)��D�i�K`�����&*��	��®�C�H��S�3��-��s�Hq�.�?�n|�lC���:����(�YQ9B�k����ԹMMc?��cş-?�������3��p-�`�����(g-[�م.de�j�S�g�X�9�����E�+nZ:_���[/׬	#{����b����<3v����ţ�1쟡����r:C!Aр}�M'�	:i�O�zQ�Z_����V7�즮h�>��M�=d�Ȗ4t{ũ�ݶ�{K/��u�h�ek�Rb��[��kZc��]���·�eo�v��$��`�$��V6����U�<�)�ޏ�/���o��X�7~����P`AYI׻�y0Գ�H�G���Osz*��2D�ܶ�F��zo����1�0� >2o�^�WO5�}���E#^f���8�L��'�����;:�U.4$a��r��m/�չ�q��o�෨1�o|�R�B" �_�L���CCvg�
�/�=[��Jj=��YD��d�<����ܼ����5�<��憱�#���C��t�>��}B}�^�;����*/3���h޷*N6����ѕ��Roh?t�PFP����"��.��r��K�@��>���;���3�[����K����h}q�A��}�?��,*!�)�ŷ|��$���kys��/�5C9r�iӫ1^�ĝ�t��������6�]��oe8�����s@[��ϻ�=)�U��8Y�~tHQn��B弧;���6�ԭ����RWR�4���m/l���z[x`�Ur�9U�q��G�� �L (��}T%�y�߻~�x}4 ���Y�b��8e�	<���^5�Y4�����ǅ��:D��'�SϢ,j�H����%E��W�O�M�4V�.�.�8��c�94��w$��+��=��ז�B�<ěz��5��QK�4i���P�Ibl�.v<��c��E��c�f˩��ԯ&
E�����	ƿ��Uq�Y��nƑ⎋�͋ �]0]~����u��(b�v���&�9��t�n��%��dp�}9��JJ�܅�4ܹ�n��+���A_�̡��Qٻc�%���A��^��93�x�R����>d�i�3t7�8"���uo� ���FY�/7�f_O��]}n�����y	X��6���������䨋�<���|�O��>���z}xV���+ ��x�z�>��e�f����;���f(�L%���7	��tT`>�YF�r�U;f�2,4�[1P��KC������y���mi�%K���|\]J���R: ���0�ӻZ�$�Ʒb��^bĎ��XO�"�^��H��n5N�_݋��-�P��*ѹ��7�W'�4��O��*zͣR��#2P�X�h<���mm�|x�j�`�%�Y�s
��<T�N�>�ݠG�u���x����W[��	M�~
f�y��Jz�ʭ����mz�����+Q��Cmv�\����j��wM�ɗG-h�3�d�a�-�!��oe<)���Ϗ�g�fkf�8� $w��:�#r��ʡ�C�-؛����#s�/�9U�#i3�����um��uc�]�ε��=��A����OG�i��a�~�{��������(J����z����4+O&�L�����[�Ѡ9�o- {X[���=�6�jO3��W2�L9��c2U�dT����ǋ�]/����K_�c~o���*��(Z0�ǜ�Ė����)�\�=� bW%��(�v�鹣�]{%�|rr����	4�')�ȼu��L4��z��xĤ�������m��O��F���c
����7� ߽98P��H`<<Gy��7��
/���b��A��񡷮��g�>Q�9�d�2yQ}y\������#���C솣x�}=�Ѫ��V8|��N��A4b�-�[�^�����A���\��/g}���^ѳèX�Cy����^��y��m�����`tl���{�M�D�S�.��Sk٣�oW����̡�鹩�Emz���y$�Ǻ�����g���J0!L�R��f׍и��خ�	0�SL���oSO^̬#ђ�+x(a����^�tm�to�d���I@l�g[)��&�_�q��;q�����=�u˯�R�M�:��Ǐ��j�y�S���ճv�	5�w����P<�m����5�mRb�s���������\�t��"���Ǖ�i��8m�z��M��y�y�W� ��-8����V����xCG��^���_|�K���Q�� �y��� ����\�_��ʾJ\����{��6V���zW)|Ȥ4�_����9)`� �:�G��?�K�@L���e9G����ڹ�N�V4�%m�.�P��i��X�D�w��^�e�5�*A�p,�N����A���dIF�y��t߂i`�@����c�3���wW�X3����-�O\o�%ͷm��9�2��?���v;�A�a�1��ߍx�\��?C��+�A��K2�U�����|�(�]R��hJ)G�4��	{s9�ݛ{P=�e��r�6k�ݵLv�Ik�떺��ͽ��p�-�����N7ڛhqυ�OG��W���1����9K�A͆�!*$�(.�]�	z��k�M��;e0J,�q����ўf�Ǐ+�l�%����k�5��6��f=����=�A��ˡ3J���=g3���U�_s�>ُUD���#N���S��u'O�v�h)<�<��݊�04��+@�\_�4Ԩ�B��F~\��^�HhDa|[6�n�^O��X��7��� �f��8`�I�^Z��LYk�1���w�7>�n���;��b+��̃�x��+���\D���,����)-�	ԭv5^��Q����h�%+��}�;]�K1��p��x~kb��]��=�H�]>���ӕ��&���g�~y���?R@��1��0��\h��XM+�	�j[+��b)t��p_z��w��x�|sW�7�W ����$��ң!�,�b�T�|��ٽ��nD�A�R��P>� ����s4X5�;OG
�=�fqڷy7AU+��_��
U�{���ȏ��{��/����q��h��6�ϧ�r�1�i�WiK�G-v�����k3\��?����3}���{q��c:�e,�Y@l�$���x�BOhF�䰼�iU�t�q�}|����.�ĭ�[��v�YNf��^���}"(*���qC=���F���;n��9m�i1�/%�LƄ],ɐ�l�a?��ͪ��{ό'�#6M��w�{�J��n!.8 �$'�܁�h_]��0�S>�2ؾ_O�����oj\E|�R�H�9���h�Rr�q�[��F���7e@�T���^�9=^��ŇS@���(Y���)�#�\pn�خ&��$/���ɶ-el'o�(��L�?�{�w� I����"����aݶ�e6?��N�I�K|�[�^�[#(뽴���7
�xM�	��d��f��q[�n�Y��}l�$�ˏ�M�t��tJ�ɧaxS��-sg���h�iZ��6?��4��?|I��W�R&�Re%_Ѣ���YCQB[O���$����']ǘ+���[� �eQ3Rt�|ڸ�E��$��1��n-�=���=���K�ٹ̕���M_'��&`�Y�%��G�R��跽(GKi6�<����s�С�"���}���ف<�������=��N;С���xNT>����ļ� ��|\Y2�G��o���6��%�̱���v$v���J�}����u��ܫ�����g�����sy��/��H�M[��* B�$_���3�i ])3y��-�����D�W��Ts6�D�9����4O��Cr�M=*tJ�/n5��ٕ���y�c2�s��%��`���>^��[m��*M�9�S����ǲ��۶x?�;�= \��G%� ~K����+�A�h-��tu�e��ǙCtӕ7����� ږ����Lď������(~?t�<�`�C%A��S��R��
�b�!T7�H��8[b}"u{g� �d�>T-6|��^}�&m�]x��hŹ nAG��l+vR�*�,�[�c����R�h�0�6ĭ����Ȏc��q�#��R�8���w��!+R��חۘ���1�{�}��d����x8���F���䑩
��ʖ�<&�Wh�������d��Z�ksS�C����rC/ǫ��G5�9d��`���՛d^����N�����u�?�v���z.�%[�����s&�R�ΟEDl�T;�P�}�D�]�*1 H��)��֢g�¡d^D����+=}g�-7���*�-�N0&I����|�ې�+ʴO��n8c����Gw���
_<���Gg�d�mq��-��>�U��F_���X1����}KI�s�f#�z�����)�D2|$)iRW���Јd��'aMaG���}}|S]�^M�Km�+:���U��'�3�&�j��{�E���_Ty�� �[Dǭ��7�n3]�ψ���r�^f��v��yoQ׎^�g���	��J��'Z���\+������^�����3?�_I�r��
�V<�����ϗZr��[���e#:AG�������=�����=_�c���]p3r[!筮�V,�ǫ��q �M`\%]8+SR#U����i� ��I�s�N�
��*�%1�CV���A�s���͖r[�Ƕ/��Xz�#@��p�x�	T����Ķ�J�dz7������ݺ�	5-9��P��%��=�)��Ϸ�	U�s#�j���}[2�w��e�g?�9w��y��������/�a3�}��R��?z 1�ⲙ��
�;�o�Lvm�DP�������y՝��f8�������R�OF�b��d��N�k���M �R�h�O��G�(��{0_nK1��ʃc��]'�:ˎ�4֋O��<�ߜP�$[�_�Ik	���)�9/�
��������O��q���x��o �KN�'e4&,[w�GbVl �TY*�u��5cF�����m���ݚ����i����ȐЩ��w&E�Gh{������v�o��'��3IRG�}T��-���<��eoi�a�XH8�8���1|���$W�dP�)�cO��I�/�����v�W)����]tH�IeU�/���~ ���#=w.���wQ�[�?:3�<l�br�� }����ʥ'�)�&�&6%%�b6����5��4/�~>�5�ݷ}nZo�Ж�V�6�N9F0E!��~�6D�|�}YG�`HX�&D���$��\<��<3DQ��U�jC�I���ړ3o>�����
%~߿��Zc�$��@��	�l�ϫ�IM�d9�y��;���	�I���:��;�ՇI����W�~����ݞY�6�W�
��j2E�/~^�A�%�#?`G[������
��O�P6>�ʐ ��Hp6l76��,^hR�u7�
��������;���Lω�~���.s�"ɓV�_�1BHP�z��ȹ]����v��)Ĥ�����E�\0r��;.oW�m�˒�b嬜�΅MA���\�;�����&��������(�W�2U@�ƿE_��j)U�-A��P��'��d���T$�����9v�c�M��N��拀ϯ�z��pk���I
���	&hI�(��Ӣ&)Xx��ă$@�.>K���Ks��]fY�A��j:�c���?�ژ%=d΃�'YKm�u�^Ȇ��`R�D�zB�ϿuB�Q�;0B�gzTa�ku∀��n��k�>f�F!��=�D�㟘P�>��&R��հ��cmLwT�od҃����o�k:9D�N��@_�����o�Ko�r�r�h��ڔ�D�-AP�M�����Z�R����)3�'Mw\i�*����7Ω�������^���l	}��.��.F|�͊kϛs]� b�g%}�6��㕟[��2l]R���+2�t���Za�s_��P#B�c�}v]�mqFAyV_�e>��H����G�ѕ��¡ɋ���Lo����h�u���J=�_�b;�~)Lt��F��/�-��URǕ���̯�s�)G�����7�D�qN�֗��]����4�R�峴�����o���׏�s2�x�#�	p�,>ЙF��2��z�h�zc�Y#�	�8)7-���^e�o+b����˃0M�'Ԏ�s���|��.��wŰ���X}Hv���	Pe�j��%/ⷬ��"�9=!��c��ǃ�>�C�/��4��[Ⱦ;����T^���C�����DXYL%��u�^��^l���P�����̻§j��zIXH��j��Wp��@��Uv����ѫ>�$=L�k7�2�vH]�
Vɟ��ξ�:i����e�7��8���;:�n젪��c4D�E��A��>\����[��>�51,�Kd��B���g�TM?�S���<��O�����?Ő�3p�D�C�Տ����6D{T�B�-]�vLa�ј��ɺ�%x�'q#5��+��)d�����\�<�_Y��� �_�>��s�����e5V/lP�y���)��ԫ��G�8�y�)��r�b��9@x���Y�c��I��97�_�����|Y\��|�!z��szW���O��;�<+�Vie������z�@�fQ��U/����1W���v�Aw��q�H�1�}�����@ d4������EUՈ�*ŷ{ceT���X�aRt1��_]NI^����>��ݡ�խ�Rqt�}�W��a�q����sV�}�C�K��=�/�����ruoƪ����yS�h�E��u�<�cr����-|�dcت�k�Ա K��/,8�\�&Hi��ō�ٴ
mN�+��k����m�6e=0���@����R�l[Z�Td���Z��q�U��*(($�Z������IWF:�Y U�tP�YW��9�* �y[�����.�*�ѩv�CJȏ�*8ƕ��r���� �7���Ȫ!�U{s��M" �G���U;�;�(���w�eTT�
j��\��)U6A�#V�4�=��w5�_��9Z��v�����_Qe�\Tk�*�*c�y`���
B��\��U}� x�_�ve��@�N֗���:+UCҁ-�
>�����K�0����Ou��ϙ����>'�P ֩���#[�J��˧8f�-��)p8��}��B�ճ����mv�j��\W���!"ۯ����kL�H�|��>}v�M�v �I�̽{�._��b�K��	)CS^Ap���\���ҌO�B`���a�c,jwr)�Ҡ����>u��t�٦� S��h3�~o����0����X�����UT�2��DR3[��'U�R�tᩗ��D�2E����H�����V�@�vXG�J�����ƥ�lc(�����⾒��-�X!��cJ�ms4GO;������Ƀ��� m���>>���@T ��R��d�CB�$�14y��������I��t���#�Kc����2��|����!�Y;��_�]��\��(�X5�lP�t�	rE�|a��A�Y˒&�ɝN��T�B��4�/1���rۤh�K����|��(�M_-��E���#`��S�x�]�x��?�v�>��9<��PdjH�_�=�A�-{>��f�F=*9˜*""j��$�i�j��xu���}�cy�zs,�	=)i� R�7����>:��ASk_�~e����v����c�(@k����b�Yy� �cP0��z�����{��*Y��jY�Ri[�x��έ��%Uݘ�
�Qօm7�G�H�����v�ܵwdg1+5�y���\����]���H��3X��1��?3�b�(���x2_i6�CR}�P�0���v��)��e{U^df�ҝ]����t�\�*sa
E�Sj�� ��<�|yEҹ` |�Ɗ"A������$@���ӈ�o2ڻ�i���%��Wq�o���/@���w�,b;�r-rB�.*��J�T%'�M�����'�k�?���73]�^�����T���c@p�F��t}�E�%%:�KM�s��1�e@�Qg�>����ҥw�J�q0���
_W�����ƹB-1�[��˃&�}�l�@L�ھ>��sTul���-kFLQQ�|F�Q�Ӆ}�!�g�i�1M�ל��mb]�~pv8 ���Wz���)���´度�Vi�.�hO1ɇ*�lWe���\$�ÑL����稔�ȣA� �Hd�-�,՟s��F� ��A�%�2+{�~"$8Q��!��wy���M>�w���5��o�#�� �6$�����r>К�
i��
�[��w��P��&j���5�r�G�8��tY��.��bQ��p���瘌�,��_��^�n
��;�x��C�-MY�c��<c�ܼ�&{���S�s5������5t'���H�����@ϔA�+������l�{�552S �W�M�ZRTЉ�oEy�:�л5W!������Tb�	V>�nϡ�Zo�{�p��;/�=�Oׯ�T����xq^+�Ų��]*h���P�����[�����H������j�����mmA��S˵�3r�%�K���][kS�3��Bm����'}���;n��ɗ��
��%�:9���B﵅�DCx� @�j��Z�VM��w�H�^#^ ���r. ���R M5+W��ӊ����X��|�w7ї +t��jȳ���>�d�9�C����H���VxQ���h<{v�k�L�)��v������qC�h8����UۄE���!���ǯ6qoK�̦��Y+Wgޑ�[S�:�LE��Nu��(n����'�����x��j��\=D5�~��A�G��Q)WA��ث�|d�� ��I�����<�o�;�9/�َ��S�u�t�{߃�m��>}�ԣk_�ii���o�1^��#�����X��b=���&l����S�<��ǧk�"EU.��qM��SL��<5B��p�zL�ҕ U4�y�#(˴#R#[��p ���c�y�G ����ְ�p}�FiJ��l���������)��0�N!��>Y=�X#�`D�{�f%�޵��&��T��J,z�-Ȫ��.c�Ȃa@9B��C�@���%1�g@!� ���6虒��tD��2�Z�5��R��BϟM�����\�X�_����Xd��NmZ5$�^�7Z-Ռ�|����ɶ��u��򼩩�ny�q/���ǃ A�|�)�V<0D�4⏾�_(!��ڣ���e5����!N�|Ѯ}K�rS�`�If �)(�ڟ)���� �!��y??+��:�a���<V��ګTS��|u�m��𶴲��{\��᢬P�g�!e;D�y��
';�������N�a%�w5��O�����X�Ţ^QQQ!���� ��h�AAW��C~t���T
 ЄD�N�Gյ������ �wD�d�dgg��>}�v �]g��.����s]�ԏ��I<�u�( �xZb�􅈂�E6�kS��.����ɹiY�I3���/�_�'�#��NE�BI�����7\����jJ�&F� ���?��\��?+�\+���~k5Z�"�D���7iZ�E[|�?/XV��g��$�L��k֗�\����j�Ѕ�S��}�t:w����?b΃+N(�������,!�O�@��H��H��wH�k�H3A'Al<~�b��Dv�t��v&�/ѣ��5��Ը�j�7(���'zٙ/@=�x�n0��ϯFKHR3#l�T���
�y9�m׮ ?�HqW{q�3Zvg�C�tXWVVFt��{�����������7Y�k#}�bc�?<�e�1Mf�''Q�ش>m�b��"��ᡡ�2���r0���D����?���J�F�Q֦1\$}���24dD�L�
M��F�ɂh��ɡ�/�B�6}�;���շD,�e��kp7�5�	����<�xc�;Dm=|ҵj���`�po��ؔX�M�f�)rx��m�`f!�5������ny��T�%>קaH�a��%�OҜ�4+�{d~��2���L}��E�S5��� �X@�$(:�;�K����W���Vw2���2�]��ܿ0(	����`B��[FRQ붳T�څƯ�V��M�=)���)�g�;	)���s�R#y�݉t�cEF��1ve�T__��(����¡\�x�d�0��y�o�2���B�H_����K����;J:Ƌ��#�!�_��*L�$��ē6@ۢ��(y&�5K�I�q8Z>��|�#$,=ճ���.+��qL,,�t�B6��|�J1��+���\��}6�9�mӝ]�����Y��W8b��b�%�$d�`�%ڋ�wc_�:������C�>�ݮw��q���m��I~�lg!m�6�-3��В�e	W.���(��� �؁D{F��D{���l��Ɏq ��%��<������V�o��?�wT�8�פ����(�#b3�Oxt���Ǩ�����w����V�����cS83Q;j:�>_��{(���8�Hh��E�����ǘ2�5�7�����?E	"��x��S�H�"@�F$8Y���|q ��L�v���=@ �n��v9�1�N�F��dM����w���{���u�0�
�Ҳ�
j��;���P�� �sD�
�**C1�W���%�W.U8��a=�Y���8)�ç����	��\\�D�+J1�t-,2����2q�?��f�Y���9�/n՗N������Kh�H����߸C"'�Z%:�����%��ג�|��$B|�!�T=����\ jF J�kl�;�nuH�@J�1�ں5(nN���z2�4��dY�������OJ .2\��i���}��&���8�Ǐ���G����;L�H��Qk��1�A�5��_B��/��Z�u6Y"l{Ox�S�&A]�ծ�E5����C&q�gV���B|XRؿ�<�+�n���M�2�i
\�0�>KY�q2T���z\�g�fm��������Yi�5 |� 9(�,%F�+W�.�����������.�ضv}է��U�W������=w�k��a���"����iQ�����:|���T�2
V|�L5�6���i�E7<������#:>�g+����![r�ɳ��>6ă*2l<;�z?� &$�� ʛ�N�9W�|�wǢG�l����S�1��X�������ؽ����R榰�
p_K�%=?�M��1<Q�:r~s�c��↹0&�1����%��XMT�Ηr)F�G��`\��9��a�9���v��׳^���j���661Ϳ���=��QX�.���g��&���|�o����-�*��o+	Y���>�f��5>PL�/��i��
�|�e��.n?���`���Ms���g���_���f�����H:�K|��Y�)�Hn�笹}:E_�e_�N�����W�C玩.��5�7l�_r����$�g�mCQ�ޱ"�ι6e����gRHR�Zw�G�e�0����WP�VD_�5���L(������-CYz��38�}����]�s���N4���P�w���|au��Ǐ���Gk�|�
>�f�`2b(�4lk��~��p3�U�gKԱ)�;^\w2���(���I��_�������&�X�Y��d͵�V#�9;^��E9�F42�̄%���Z�+�/�9�KD��=n��0S�eՐc�98��bvS�g��.���3�&)U	�� ���)4+�4RMl``�ғ&�f�;�H����8���!�i�����B���E�,���y�}���y�6,��ųp��<[�H�-͵�ʾ��K��,vĐp�q�b�0Zn�k��p��=�5�w���!BO �d��fF���Pj5p=
	>JX�Ж]�ƊP2���i�E�rs���� ��$�4�ÅR��,���te�Z�@N�E=�}�6�e�ࡋ�FD�5�ܹ��0T��R�7�&J�2�m8�|��m�s[����
G�{Zi4��j�E^4��S744L�	C��n�fj��WL���\~�Ր��Oh2��@v ������[nWI	_�6�x��ּ�&0��Y�)��'�%>�t�Cm&R^;��a��~_{�DHL�#��}G(���ľg��	���ZL�d�l�+c���d�	i�,��W���g ��Y�/�2���ԗ�_���8ޑ��0ś�C丂��YzYCG.~~����\-�*$HD����Hq�^ � \bd� ��D��EL�qq��<�X ��x��	�`�i`��Ps�B�݌3����_A����!·C�i���ie��K&M��Y+F�$�1LYL�OnPP\)k��KG'�\j�J���R!��v�'fk�r���������8�4m����eVE�^ջlU���7"N��]|���}�Qc��"W�zpYtu(?ߙ��9�!�Jۈ Е�>P���#K|�D�ԒE�#}a��k��45G��`�A�F�����N�xS��k��[J�ٜ/�י�y��8���,�Y��G?bG*_��=��&>{V�1:��S���HG������djc�k�@��u3��եO#o�ҤW���.��~33���n�G��?�a��p����u�G�Qc�� jgA��$*�s?^5�Y����Z.2ͻ*)�K��ƹ ɗ��eQ {>�K�׆g��ֿ??�GH��/^��D��T _�2���ױ�q#��'=1p�$4@�
n}}��P��=��`��a��aF�(~�j�~���q��
>[�vݞXOSn5�N��=-+ݣ����ȺMMh�T��j�����^�"�>��|v�����$�oc��Ç�r��O����	�J�_`���Kz5��hSX��ŝED���d�"������Jry0u���&����b��Y��.ko��R��/��n��+r[#�r$!��;KDT��zD�|��*��I¬���#��a{ؙK��cb��^1��v��u�T	E��_� ��y' �[~�������%��=j���r\sJ��e}W��I�Ӊ�xB�
�b='���8�3�7É��}���N�7�{��עn̹��:���jAT,
N��.�T�N+3��Np#�N�a�hВ�R7�@��� ��I[�sJ�"��Y�A��"J�z>	���e��ྐྵ�g�2�ۯ���K�V���Ԃ�C�9i�[�*�}��Ar!n*r�A�,/��"�C�U-{;=�������մ��ܻ�M"�~�񺻏%��
�V��j����]7�m�ט�|�#�7�ѣ�����zZ�C�U�z~�Pk �z\ ���~����&����;v��	�j�ޡ�\&cOZcp�Q��G��omq_���Z���)1�He��Ɋ��Li䘏#\�iN���gpΫs�K����=�ob .���F+���iw5���u������E�ls�کz8������M��q����㶧�^�'{����5[Ēǻ}t�������,��ݟ�B=��Ѓs����~�����=����n-o�'�5@z	Q$/Rj�Z���ݗՌ�-+j����Z�#��E0;�ǯ�8�8X�k���ͷ���s~`���`g�O>�i!���t�Ld#\h��� :���g[eZ�Ӭ�d�q'_������p8|���h�|ߥFH��	΍���x�����hD���FlHHH�QS`o���󡢋��k���&���~ӕ��=^���E�����|�v{�i�BhG��v_v�r��̢���Py&`a�Z�w4���~}��h���-C+?{'G�u9��g�����$������kh��%>��Q:|��7k��$�^��� C�[�n���jݫN+��$ �5N�.�j˙�߳ԛb�������v�W\BO����S��ɮ  ���԰�����N��[(�/ �[!�w|������_`{���M��r��b�G*KK������4=���p�1,G���nwު�D���>��Q/.##�ߔ�[�w�+��.O��|ΜK$��6vB�j�b�
���=b���r���,+��4��M�?Ca�8���h'9�u��Ap���_{%d�+akl��]K���PP M�屐�z{����>����[y�T�,��(a�����q�������8��)�0���(��T�yj���x>�h>:"�k>�.�5x=��f����S�C��7 A��F�I5Z�#Ƒ�Ѵ@��9PT�'������[=f�3���b8"��&��	k���l�,��F�,6x��1���|T}��}���Y99�*�V[���F5W0���c�݁���4��̂w�di�n=Y��59l�\q�j�:Ͻ�����
�A�L�L@�#�H�X�`՚��$5��7��qp+��@���?��rrr;��TN���A ۋڔ��̝#��[o8�?2
��%���wZH���jd+�'v�;L(���K��*?	������Uy��YrՉx~�&�dK|g�4��n1��y�m�P0����u�1�(�Uo�U2��up0�χ�s�{�G�(�h_�U���;cBٞ�) ;7[�|ݗ���ʔ�~0���u����W
�E�� ���N�$�= G�1��i@8$:ܕ.��^�r��:/��V�(>�z�ݷ��	ʥ�<����������s�l����8?XL�o�����;�E��19��t�����&�m5�p֢��!خ�T]Q����͇/���<��yR7�-r�G�6V�ٛ�!+V���J��JJ�ۑ�!�y�Ȭ�-�F v���2H��t{W���RK>��>�7� ��]IT�����A�;�pbE{�A��C���kd��D=����^�7.�~>����`������1�Y�����K��yS"�婢F�KRP p��m��>����;ٿl����T�y�Zf���"�Qw+Row�"�*�'�cp�"@.��J������i���V
U)�4��%���goq�Y}��g��b��_K�$ʡ"��犆�WU���#��)�?lL�+{���i?Qr4U,��|B��n��	^�xe��_l
��S@o�H� :���f9��M�D<�8�!�$5�%%�2ہZ���FF�oĢW^Y�%���y�(�x?�|�[1��u!� �I�|��ˤ���5�z)9ɣ}�t}£>T�I@O	C�ek��������V��Zf��F�0#��!��@k�HEQD�Ϫ�߰�!��c�c��}��3)1��H!
"���0��AI� ���H� Rb�"!� ����tw�t=�0��|���|���D��}v�����9�}k�>�{f�}1x��L�y3��]�W8Hr�w%<%I�u���ş�<�\�^�M�ܞ�`1��G�ɇ�-]r�-#(4s��؋��h�!�+l5��/k�OG)�y�;:��Y���Z���!FYeeQ{�*��ɩ�޻}�q��Aq�M��L�W��f�F�ISW�~p^V34L,8G
������h<Ay~�1�*���m��Kq�(MN�
p3"f#�eY�;*�������l�vk��ˍ[��U��Hv�P0�*�O�Ư~��uy|zG�P���F3m/�����f9�<�'��/�"�٨F�8څD}�D������R��@�[.l�AD��u��ʌkV9���՝_ۓ�y5[�Ҩ�� S��	I��S������桸�J�)�}��5����B�6F�?���2Z�*sRIFm53&V�*���V�IW.�����(�Ǆ����P���z鋱�R����(%u��p��8@�^8E�?��ti�k�T�[�0�W�Bb�F"�R.+g"_��w;�f��XTO4��YB�/&(^�<��q�#��G����?~�e����չ=7B3~��t�	�6�	�>�i���8�ؽ���{+|Q�1
Ԩzl�ύ
�$\�9���֬ᐈ��|[G��@M9�4�!�#� m#�BKw_�F��H�
����r�Ӌ_b_�e��e4�J���[j�8Ze?*2�V�pL�04��W���idE�mN���y���n��m�g�������*����y�-Lа+�E~6t�Y��R�H�q�U��o���c����Y�1���#�;w�y8:)��ο�L8~��[<���i�l>���Ю۳���#�G)�Ч�X�5�s��SM&�������Nǈ�.P�� ���%�׃�+�t���ߤ���R�`�pB~�8Z�O�H��Y�Ό(��(��@/��q�}�Y��=�����G?M��EBE.Mmm�[����y/��l�KNo�HMn��-�eK���h�~��F�V�ş��V���y�!o4����㼚��O
��?���-g}���M,��L0�X���K ] ��,���MBdE#�	��H��̆mU����P�c±|����sJj��B�'�0/{���d�pY$��󌹺��[�5P��";�j�����k]�>��z_����M���Z���7��A�#L��\���Z���+�����5D� ��`�+�t�,���Vx�# ��Mg��n�l�/<ג+�C�}ӶIv�F/�Ä(X����4���)ϔQ�e��}���˗4\����U�i �̚Ż/�,ƻ��[vs㟎KR0�儚2��!H��Q��H�r[���!���zd����sWlw��ϛ��ʦ^�}G33��� rQ��]��/�J��w�Ѓ�V�k���7��o�z�lq�_�2;�� �OV���M&������T <d���M7��iܥ�Qγl���'��5q�V�zr&�^���
��FZV�G.b;����4����l�u�ȎI��Ω�C���ᑷf�:����u�4�a�����o�Ez=QD"���~(�k������
�$UՕ4�$kjdD�ȃf��]� j����/"`��G5R�u����7w�`i��{���]E>M����m3n����1acjn��Y���ΰh��6�f7^ACJ�Z۝�W�U�:��S+���gш��u99߂7��@�S��d
�l#��f@�o5�>����8(!4��^�h��#�& ?/s�ӥhg���)W9�8	�*9XKn���/�sq�>�m���#��G�.��}�%�f �w�i��J�����[2�|���Օ7&��!t���PO=�t~�8�����c�u�6x�\n?)�M�zU�8Y�]��573���ڛ��b~���������Kp�/fw�_�acɴ�%Cyw�q���,��r^������H�|A	Q"�4�7��`ɐf��Z[gƱ��ܳ&����~��Ss�1��D�q �`q>Nv�}<�k2���k�K�d�����(�,N����P�Lt���P@*�S
�Ҍ���ßx�V��`9/.��@�����NBA��ZU_��[��L����M����)5կ�ÏLw�Z�z&�,Y&ǐMl��6��ÄQ8J��u�r2ء��)B��!a��r��Kh**�	Ɣk�؞�B{ňXe�8,���_����ܟ�d�Wl4��~k��S�(؋�@q�]�s���v���>R�X%I���#oK���������i��D�q3��wnc~3m ӓ�'�^�T֑������nn)z��Ռ��
���'v�I�I�=�{*ֳ��9��Ok�8���D~5 �}���x�S
[��~.�V�"�Ö-AJ���n��|��mP{�X3��g�����f��M$�pp��s��XnIe}���-��d� �Xr�92��,E�D#ihE�� ��Vn���|f��h�%���UX�c`�z����(!NI�/;N������:=���DĖ��uHΟ�@j��:w��)ֵ�p�I�����0^z'{��՗�ϩ����u_�ׇ���;A-a���%Z�۠?�#qg�4�:�+'8�5��m�%G�b�W����!l��Ŷ2Lj�G�r�}cp��P��{�Q�b@>�y���9��v[���B�����{J:�89��4��0�}�N���h���k�h��pf�\��w�zD��y�:�.ǎ���Eԧ��\� +��m��<���e2�4^��ٴ�A�=f�	����w�m��B��&2	��4��QbF�:�[���w��9N$�G�	<��ARIQ)� ��^(|타!+�_�ڹ(	0�rhR����Zź�f�y_��Βl�^�We崨�Kk���l�v?z��}ͯZ�S�g��y��пg޵L����L-.fۑ���M�J��r���jڨ|�X)!_���Fq�1KXS�Q�,º��)����Ge=�C��_���t澗���-�2V�R �3E1�1��ϡ)
b�Wr�c�����
�i�?�	Aߌ�~4�yB`�n�R�mW����3�\K���b�_���}S���)f�V���q�"A'=9���#=2��
����@o��$(��L��Ʈ���~ҭ/�<ww��FG����so>�f�6+E�pS?��;I��R��F�׏8���y7�1��M��	<����N814�����J�rvۆ�����W[Yn۟��jbo�R0U�Ɉ�
����Ρ<%r̢��b�"�<y����˗�=�Wӿ�4���Uh�ob�rٚ��R�q�����}˜��6�	�t�U��ڶ�F�,_a!�X4����bL�^)nxyOƃ�Þ�"^���=7���Cv\� �\~.?b7#���x5/oRc�ʭ�yJ����6u�}�v��9���Fsk�B��ͽ��j�+�K�m;B+�z���Y6�]�NUs!0��]�<�qȓ����<��I}��b�p�/d�_��Y<eй��W��8�j��i��K��u�O7��>�0j�oʓ+n�~�����߽GyK����/�B_���.nJh����Ta9���G�P� a�A¬��enN�����o�(677w?V�GsX4d=BM���o�S���[���X�rb�}�p�ö~��M'4�+��Ÿjd�\p�c���}���6�-%�?\�և������7-��I�X4�T�I#�/_�~	A�����=�(D����|�,$E���]Al<�����N�i��έ�ƤGi�kl�'����9E��޹ل,����s3�6�� k�[�֬j�dacs�@{P��[�����t���û�ڙh7�'�l�b>ɥ�+/���Yj�:d���?Mx�q1�۳g(��1���k��/j�y@J��3��8� h��լ! #��v�n�I���ec[��v3�L�pXr}��Xt�D�	����]Q�p�_SI�nD�௕k�9,5�__����ͯ��d<�O�~�|2\�9VzHˆ���N��n��`��4:�-y[��m�&�(nc�4��騄�<on��Y��&4�m���y��pz�e�$�۷���KD776��su�:��d8F�$(-=�ֺ�RK'Vdt��k��Dq^_��'�0�����RM(79(q��Ά�m-�.6�H�5``,�E���� �2��|�p��O��''}r�	n��_����r_n�ʦ�~���~�eJ�奞��]��Lu�斖���i�P�b��(`�sl�����t	l�����:9B�Σ��X0A�	�>A�%_��;m}��\B"��� �0���1������1�	
nߞ2��Ҹ�o<�P�~T�'�"��h��{{6��l*�`-/T�q�����'����.��6��嗌�?7L:CxF��X�H�?"*��ET%�2z�w���&�L+��P�Q���%| 2��i��AQb)aG�.�4���pǞ�� Z]��r"��1V���E�2s�Wшd�?�O��3����f���7��Fu`F�=��J/�$�
س�y�&�OT;�?C�]��ڌ'���;�~#{������s�'�6�b���XS���%fq�d�b�!����,�1q��.��+�Ÿm	����8�~����؛��`͊�7��%�"=�K�]�������%?_�s���w��炧�Q k���W����>#����
��T�c�p��B�8���/$X{�o?�+Ĝ���!��Ē O�o�	��?�I�VyH�##��nJ�(<q�o�y�!q
/�O~��_�[���MAS�>o{�3��D�-�`�r�V�6����4�7�'nx��[��.0�����_��M| =�[��(mY?�k�(��$7���|/B�j�(�<cD��aHd�hl����;A��>s=tN��w١ˢ�������L�1��j��G��c���15�i{H�I�fǙn�����B��7
6"�Щ��ؕ����w/j�8>��4�a�{n�^;�+{���^����S��d˘���-�LS��W��jtj}z����Gj4�!��gN���U,�P�h��끁�#����,����-`w(e)|w�1-��&s�K�T�^��>�/U'�8���o��U �fax�}�\<�`���p�F��z��92�����m)Jj��)���)�^��	N6�A��zh�ĸJ�\��3~�ß�U�ylӿ�a:�4�N!a�Jd[�P+�}*������b=_�A2�\�Gr�Oe1DD����wB�*����� �����^�J~����1SԼ��J����U���L�7�5�S�~�����eq_��>�iw�,��2/�ϟ��� ��2~A����ʵK��Y����(��|��K�s-JEO��
\�����L��~o�[e�륰�����Ģ]l���i�nZ�?�6S7�|`�
���4��:����(Ő!�ݧ��\������6��߁��8��Bl�f�IЂF��@�dH��;����f�Ը�Ƭ��V�x!��v&'7wvh�3��6�^����m�^�d_� ��3YǼr����%�Ȉn�����s���Z��į��[���p�IJ�װ *`�Z{x1��/�HC�f�������?z������m1�~4�8��
<�����@ܞ��B��ƺ�^2��ѷAEs������7��QoG�	�I���>�d��)j3���*	Rq��33�K�D�Q�>����!'�+�S��]16�[�u���O@��h�i3���T-�%:Nx!n���*�YŌ��S���=x���_��o��G���sw~{�����>`dG���]���_�R��x�z
S|xyJ[!R=T��-�<�~>�F3�s��Q2h��T�r����f�v	Y��8|\T���b웸�ccg���͐������}�3N����g�����$�3������r����	�L��J�m����W?>�@d)>'h)�u��I'��.�oeh(ЏJf}��p�<�� 8��B���b�
K���H�"+�?o�,͆S�� m�~��o�k�޿�3*^�~}[eǜ�;���_t*�aM�s��^�����,�����U�5�W��/7���Ko�p��&���ō\��У2t� �f��n�^�{!��]�-���'5n�/k���kj�K�������S����R�{!�#�ڬ0�o�UlzD�P�4�&����`�l��auT�k��d}=��i�"Z%=��Qہޘ�Da�a��g�ڞ4?t���b��{z���R���1O0F��gW����ܻ>�=��ш�~�t!�]s�M����8�����G�A�}o��R���L�bRZ��c�?f�F���<|��m��0E�ܜ��w��˩�=�Fl %��.
ըHɬ�AӍ=����m�X%_�H�Nˡ�����������▊l�tSb9$+%%��qGۃ0俻�B�./O���mF�Z�~������4�ϴ�OT�<�B�Q�mP=�0��O4	��<Zޯl��rf�J!����?H%���~�/D������o�܋��_��e���	!z�`T�5�j5R��gè�l�v���XDD�{<�#c%r3���+�o}����mĻ+Ƴ3��r�͉���{�7����bv�'|�&�Wt��r͜An���<�8񢰹Zq�p/X�?[(P��r./��r̻�����.C��1ۋl�9v�jd;fQ��=)��?�-7���;m������uƧ��h6�H�I�y�<i�ki����.����jx��G��Z����T��U�x���>H:����	�j{e�v��e��Ňw�L�b��!Dg���������H_��?k��Z��j�ְ�v�h�8H�N����ρNq��e���<�Ҍ�*��4�/]�q�COQ�'������I���#�%_�3��=�Lz��\�o�6������)��΢��
� ������IF7���E�󬟛uv�&G�����_D	lA���S�{��?0�����d:�	%>�"�"��pDO�K^+�u�y�c}�)��R����'�������u�s��2%��5�NSqU��>��O"h��,�܎t]u�>��I�`s��LMG�R�ʧ+�ם�Y��:�1���w��ݎJxG�od�o����9d��_�*wE芧��Z�6T��i
�>n_r�� Vb��
����(чC�Ŋ,��nM�O�Fb��r���y�\$$�V"��v��A�p��@�YZ�O��� R�Q�P�u��L�GxO';::�<ĳ���{�ꉈb�K�X�����+�L�����/�h0�B_�G�%��F�{��@ �d�i���ǃ_�W��\VO�������o�Z�'��
���.30^��-�9;[��B�R:#���'EOx-��W�Ŧ�� ��W`KK(��M�����~�Q�� y�+E��}[^�Jc�#�2kmW�툮%_u�af})�/�!2	��r�ч	Ų����ӯ	*!;b�L,�SG����6��]�-�} �$�������pv��ĐP�K���NC?�^�@�`p>��k�(o��fF%�2>>�W��/�O��C�ӟJ�%�P�+aJ�l��+Z�����\�*��6�+b�?����;�-�8��|��F/�+#��4�^03�e���j(/��ړ���I�����;��S��JO����"fS��
K�+-�{��|=vb�\�f�+����"�v��1�$�.�	���5U*���YȎA��j�����7�e+|��X����I�@���6�=��׻�ggʞu5-�-�'W,8�n�P,�I8�7ߘl�-�"ד�ԽoU_hw�u���ޙx~*�+�}ǋ�r�>�qF�=��͞ohS@��g���/�0ǳ���Ӊ��_jI����+X�����V����M��8$�7�쳶���f�9��h
�EĒ�Q#���^o��Y��R���mGΣ�E�xn���T������Vnp�VE���j�Șō�!���kN?%�"$T_�/�q�-$k_s�wx�{ē_)�.��a�A��@��X��O��B�Щ����M�=�|VQ�f��:������g%��K?l�X&�8�O�U�^�Y���Ý*��\Enʕ���G����@x]�>�3�ӷ���pW���#���T��և���lF��Ŝ�^=ng�fm	4L��]�rV��$f}��=6��,w�K�����h�[�J���O�kL����s�T�l�Z��Mh��f2K�[M�� J���$B�*��p�R�5�2���Z�X�(/A�U���Ϲ�'L��x�p�[�
����Q�XL��o�;m��%*?0DX{7>B�w[k�h���g}�����i�'l���v�
*�Jw~|�����Q�]G�΁�ڥa�9�GvQ��]4aZ3柂jx��?�Y��dP��D��U�#������x��D� �A��&Hц鴋s���a�:-���:i9��T�ų`��j3x-���p�� 	�����n�>����[�j���,8�H���/T��{xa��W��8�Y1�_Xì�k�w�����gØ����	�v/1.b��\o���@�ܼ��yx­0ЅU6�r�&O�`t�Z�d��2�ź���,�:��߫��n?��ʵ���B��G��Y�  CTQD bP�����%֖�`�֟1k�`
�cPfaVF�����- �:�s}����>Z�5��Fy�	F:�r����X�{D��-e)�W���f�E�zf�����l�GS�^h.�x�.[N�ۓvHh=��V'��Wd��v��^7�䤟z��cE�A����_B��;���l�}!ĉa.���5�uu.�Q�ի|a���u�R���i�C�}����4ŉ�=y��>�����S� 0���P���tFe�a��_Uk�|�?Q־���_5C���Wk�ԭ~֡�LȠ�J�fDE]��!�n�� �� �
���I{���n�靨*	J7�s��ܷ��E�%�r�k�o��� b��q"��7�\n��ﲇ���o�[>��㪀�B(�������"ڴ�%�(�9��p�Ih��4���-��[~q\��\mt� y�S��<�k����W��GJo����㱚L*��^� �J�,�\�X�!S#.@&�J���,a�R>Z���8�����Uܳ�\�N}���X�+j�'��Тmj�:��fR�8��_?���|;7ߒM�_����4�P�zP�ۑ+9w��MK�ݯ�@��B<.�A?��"An�	�@�jH��^[��y���A���!s��3��d�퓱H�ş������]�Ǿ��yҽѕ�����&�5]�>�����r[0\s����\���~C�X�'qLW��$L^��t�O�Cc�/�����KƉ{�~��#$!ѥ�!Rvk�?	ۆn��h���y'�<(�/Z^^Wj���I�#�n �}O�?���<���:�U��88�{�&AR�t��Ŕ���k����'���9-�W �BL��![p�i�Iآ�ݡaM����lKw���H�����c>��&�k;Bx���*�o
����C5u�u���Vo*߽s{��u�d˽VQI_Gϼ� Q�z�ˢ��F�m���b��,��V���<}���˙�h#K4��P��,���@�^$�GI<�qg����-�4C8��{m'���~��p�lt�|EI��_��>QL`���-��g�-�(�:h{�(!\��_*|�!������RL�J�x�����kL��s���T0,�q��N�p�V�7�u��yp;_��k�FФ�ݓ�?9�'��nC�EEį�����*k�2U�Bz��fk�����/��N%�ZR֜P���`��[J��A�4S��s����~0��l�6@���B�9���zl8J��[�I�@و̽`����������m��q�;�3�ۏ�u�hҤ�8�z��۾�}]"y��$�Y%ӌ���p�B��CMٻ�C~��^�8���������1��B�pg~Se�O$%��ޯ/|�v�4S�DF��7(=����3���l?�6N����m/t�r�����_�x��N�J�|e񆥏�>^���ڗ�O���h#UiT]��`�)U��v��իq�f�S��ï�P�n
l�R�=�b��r�w�`�`�Z�#��
 ��g�ޢ��Tm6��h68�qӄ�J�Y����{���fk�f�I��Y��.ϳ �K�L~���/yW$+��L�
N��k��ެ�ϝ��t�6��^���/�{��GQ�Z�&�}�� L��tK�ꃱu�����,i\�uI5Z9Ha[����p����egN\yA�f��J��[
���~�F���qO)��Ӎ�'�qwY��n){F�j�b�[U�Զz�������l�����},�RU*�5���Ӑ�cYՉ8=j>�Db��k�s�"s��w���`lc�b-D*�sr��ӅJ�>�����@��Bȫ��~�p�k���[D�b����;�J5��x�q*�vx���}����TP�j����:�/�Zys�w�AH��W���\\J�ĳ�٧�xJ�yE�A^��?��ӗ�5�g��w�١G����^�V�;{ǔ*O#;�\����ߢ;^u��l��a`J���9�7m�@(�7�=I-�Ӈ�<تP� t���{	`1� ϭ51�8U��xˤ(v�_q�8Mw���{�⛭Tvg��G%yL�hOc��j~y��J`i��éqZ)W�89d�tj���ϟ�/*l���.
\��y�eMAA���_�=�ҽ,�v"��ζH $@A��/J�҅���n_�$��"gf�%$q����Mu��f \���=7|1ܭ_�,��:'0��r�qS*�Z�XTd5"���QFL7g���}1��S���h<��$�p���<2{�<l�~��st�Z��h�_~��)�3xK�8�N��@q�?��Xt60T�^�U���c������W�mæW���9�s��䌮פɼ��L�$�eĻ6s(*��A23�M"�~�A(�����7�l"����-�:\��s;��54�p7f���˗�Q޶4��5��"���d)zQ �������0������]��G�?a�b����s�b7\??,����oS��5Ԅ�Zw��4*��|�"O�q���;8�5(�/��ٷ�*++k6���[�,L�k�,�uzQQ$�j��;ojCRFr���ۃ�}�;.�����5~<,(�t��9�۷Ix�+ܣo�/7�8_�@QƈX���҇v��[�5���(�N�]V)�HjN�|� ���KO��z��Ï��W�L~>,|�+�R$�ϯ�53f��ſ��=*����	^�������|�y�G���V:w�^`knnI�������=Ǎ�J� iX����.�\�W��5��X���sc:���J7��ӝ��Ԧ�&w��tb�bW���J�*H �3��N��i{��G�x���ub��Tj���={ ����M��f<\�?���I��mV�I�%o5����?4��O��$E�9��_=�_x>��>����çrD,��꺆����օ�Q�Xm3���8	m�v}��6� A?�Z��S�)��,�?��	�7�祾�u�`V�E_�u��BDn�z��3�����ӄzB�O\�С6�?��	�n��E��L^ǐ��NKE�zw]�_���&��#^��=���i�{��(��!6�h~�՝����ة[-5C�%r��ĊOu�|�����XL2d4��U`���Z�o5t��̤H�I2�9�R��ؽ��ء�/Ӆ.`��yi��C�)�;L��d�H���� ��g[)ie%Y"����}<BO��[j`����4I� k��qVG��/-�������T�h�pR33�6c�3��#HךQ0#W?@��ӛW�e�V�G��bY�jL�u�`����g[a �����tu�Vʇ�솠z���s�H�@�ԭ�p}�e@o՛�z���~|z՟�; �>��Y�2���I�"�?�Wj�]ӗ+]e��]�7�s`��i�OId��8�HF��I�FƥF���+o�W���ϝw�[�����]5�~��ُ�?�"����w��W�W��X�A#=�ǝB��4�TxH�ܜ��t�l��GIz|kvu%g�Ą�! �Lg�����:�#����I������֮�oZz~ŷ�B�������b���&�W�1Q#�R��S�ZɊ�~��J�w���{��P�x_�� �y.击�V�_K��o��J�9s��?�j������ȓ�zָ,G9���@�̘�>v��[�	S�F�, �wGg��G�D�ݏW�T����2�Џ%����G��;��mf���Q?c��p���Z�n�#���F+!�L<ÏH2I7�d�㚠r؝'�I�<M3&�Г�_�&��X�o+2�ǘy�Q�V�ͷo�WdF,�Vh��v��Mft�'����,v'���2�o]���{�:��Fg��m�5u^�7���rq�wg���#E���=Qf�]��f#y9�g�����.�+g���A�����b�a��gyX7*p:�<�t��:`e ��F�} %̺?3lo��u{�z�C�,G��k�G%����R��_n�F ;�a��F^$��Ü��,'{s4!7Ĝ�v��R�?#}��������������TX%��κ�EgOB5FY�~H!ru��_����+`���N',�@V�m]630&l9��їo �$`��Y[�^ͳ��A���������&$��������v3��_k#�\�_$����En��ϫ���1�>�Gx�Z��<���j<��\���O���;������P��0
�.`{��NT����4Q���m�����Uz�/�#�D��n5����3Y=�R5|,4Vm�`K�+���N!�b��.����gӀl�᜜�V�FmJ�Gqeۯ7�	n�}*�_�ig�?'���b�߷�rOIM���6����L�x����٫s�y�'��]�bOL��@W��3q����)�"g�w�3a��ݭU�ݾ���tϻ�b |�iT���Z�/��e,��Ȋ���R�~G��\����&q��3eO|�v���Pi�Z���gB�h��tN���0أo��뫟�>��)8���.��p�jQW�8m���Q�S������o�;ˠ'����NK�?d����O-sMdV�sĲ���GQ_���B`WVjHvL��sӾ��{U[�1�%N#���~�����Xx��[�H߄h��o�M��2O'U]��x}/�~�>#^�P�XH=��P���<�T�][0��l;�:�������VtNu����s�̼�^aѰ�y.b�mT:]O�Z��T�ܵ���t��(.���F���Nh�A%��Ȓ>�}� WJ�郔�p%>q�U	�2=U2LRL�!�$4���`e Ng{J�O1�,�Q,2cR�ӳ�w+���ikaҌ��<bs��k�e����H���V}�{�3�u�.$�0��2�f&p�.\y�$,��cE��T��Z-\������,��~�"�Y�x��tR�j��p�t��e^xu������Ւ`��R���3�n��g	B:����tMx����#��l῰����,�����D��<MN��ݲ����N>4`ē��@��,m�b��p�\��'���E���Rϱ-�p �2�3���r5�qE@�@@�Ê��!�~��lq��<Ȣ���b|�̓W{�P7�d�&��j��u��5١�I��e����Cx����!�g]���p�%��0%� ����k�����]Qb����)�_pPx�"�1f[ٸd�@,&�}���e;���O�q����{Q<<u~2�P�X�h��eЩ^=�c�}B�Z.z�R�Cw�5,ߨi�#��PH	���&�|H~�/*�Kޗ�~�����.6z�������--)����{x���l��%	�"�"����:rr�MI���G�,\2��������ZzfHf<ܭ�麳���$p�:筨b�3,R[P_�:5�w�;9�=,&&�����Tg�)�'$Ʃ� Wp��喎_���j� ���ϜE�B�r��@�p>�ES��W�ƌ�4"�m_���G�#$5o�%�L�w�sg����r��;�� �����YL^O���bl������b%�v{����6�J~�k��<���x;�o��%�}�/�q���.�r��'�Q����L�T��bl�����/���)_�9MB�ډ�Ę$;�//�~	�U�.�譞"F|��N4�u�+%�!2�N�m$zh�ǳ���j}W99�.�<�H���<���J���d��>���@ �j�J$�g+�7�:���p	�H��/q:'&	����Nt�;��-���'�ݻ�ݿm�K�"p������ϲr������7�g'��� ��p3ߎ�yQ�k:����%���`�Y�ED�c�=	�zo^��d��H�����O9X9=���2-��k�JE����y���-j1R�E(�ӣ;i����扊	<T�a�@O��susu�E��ƿ#�\�����&{X�5�MJ5x�9�<?��D��\ �_����^�`?��	dE*��� P�z6#���Y]�YX�<��a��x�kt�����O��ng�����G	�$��2G�4c���s�i{�+�J�u�Ï���u��С�X2S�q��W��~.q>!�
�� /0[���tM�x��_���q�oo/�p� �q����\�g}��ۘ������# %��4U��#��uƦ��ѡ֭��҉BP9�}r��߿㪻ro�+%@�s>Hb-��4X������{��9�	@��̋RI��C�?�M;N"�#�Xq�3�]���T�vVa��a������?�Ӫ����O����	���_���ׯrx��k�X񒳏3�ŵ���kO�����(�:��3�1y ��/��	
�(E�eh�ȗ �tzJ-��,5%c�. �^�pHF�TN�����^�`?{�6�RK�e�%z�۲))�4��t�����L�v��r~���$рa�"��(���J��ad����Z����8g���}�/�'�^�?�C��o��x:(J����	��WE���Jf:�����~�~~�L����Wy*���\�z�������H1MCK�;,�þt�@�/5��h��-��_�M�\����z��Q��3_�gM���щ9ñ���\F��uM]��(�h���I��2��TS��s짿ӄ�6�>����kn��w7��$�4ܰ���Q��7jaMrO�>�P3�E�4������:��P�2OE �I�� �01*��pe�$�6�趹�y闑�J1��Q����h���MMM�ӣ=����.a�Ӄ�"؝�*��i4~$��������s_M�u)
h�N�ȍ�z�z8�??�C��pSFj�k�5=�c��Co�T�x!N��Ύ����������֑?bۉ`�t������ڒ0��.3�;�\�E�Ue��@�u���d��!E��tpe�ܦL�-�+�
�ќG�����@S;�('b�8��n
�������3�eq|�D!�0�Bd��=��+�4����2?����ŝ����E/���>��ys��Y�kʽ��K<� �l�tV�}~���@�A|�i�U��SAj���g�e�n'�ۭw��=P���r�Z���1��{�>�� ���ؼ#!_��.z���`x��ˏ������o��|�a�^1��n�k8a����CG�\�3;��nh�ū�ؤ���0�2�;�njU�X����!M�0������!>�8. ��ڎ���$9=N�š����;��4r�4}�'b�����K��zŻu5��U�]xuwT�K	U[Bm떐j���+I�ˤ���\��<o������<t���V� d*���F^�l�}�ai��*CgU�Y�����ާ�xj���60���[0�OZ��m�+uz[�3>R�5����ۆh2��z���[z~q��Qv,�.��kh��,:B�8�t��@��s�J=�p@��o�g�x�y�	=�t��2�<�]IT��T�+hŶ������]hj$�9i�����O[s��y�I����_a�v����&�_�߽��9>���{�j�3&�QY��@�'�}���t�ފחs'_�׮�ǾU��������6�N6G��#V��2��9�d��@�_��
����,��a���UBey�.���\�6\c�$��{'�}?�kE���>��T5����c�v� ����f���Qi�������z��Y�����K��e��ǌ���Tyg ^Aa��&�G#�o��}�����I�Җ���DW�n�v9�wJ�COs��\�*O@���:ͣ&�XJ�?l:=��&l�Q��:6����ut�>�?0�[��ӽ����oö���E���FZ*te�����aK;�~���?Xh�ۤ�7��}�{:0��T��a��C�2!���F)v[�]xo��)���r���0���x���]gq��b2�q�ՍI&��8N�~���pT�����eD�N�ưLa��M�6�X�R��	�Qڬ�R0n�і-�-�o��:Wx��ϱ�Q*�w�-�v���m�5��mD�9,R�i��p��^���W����m[���oE����������f��	�1�r�V��ű�>���Z�U�+fff_^����\J�]�/lS���_�<�D��5M�.4jx���˹O/-¸[ch�D���Sg~U�v�M!��[�`���t�v�����\�r�h��Ks
�*�4�Gz���v��k8�M������R��o][F!�A�/���_ՠ淣S���z���⏨������vN��ZE��ߪ+�8
J�R.�b��p��� ps[����_���A\24C�'�恾����K�y���ZLB����`��ׯ#�%%?�u?�K���O���\���~�
ÙE��RN��ç����n�0�y>sƐ�N17@�]4 `\���R̜�҃���Zfc�u/���vSJZ��o\>N!NۗH��W��|Ʈc�������3M/��m�<� $:���'8쎊��$����ť���~z�!��Ʈ�Ν�e���Nz�̿@��Irh��c#���`M�x�&� {�������J� �=f&��ܶ|}}�R�
�=�(֣�҇�xD� �}���z�jx��xN\rt�d�������zh���ܾ"nJ�u�]��v�B��아��5��]d^+�Y�w����3��������������99������x<�Ko@o�%դ��Ǟ��R�Gs_wI��$X`6g�-�ǿ�D�$����{]�z7-X��L���pJ�{r��[��#�O�W5��S�G�R��8� U��72���	9���f���3/2s�k��PU�!�j�ǯCO�_'�w�2��-g�٘L4<��wsi|����ؒryTe�퀷�1��Ш��Dtp�<W��(��������Z��p�ଙ��׳]=,����]̙70�[/�!^��^��C�,^�٬:;>{v��:!;��5��`�xǋ<F.�1ZSgv0���u����Ն|��L� ����Q���*�>8�^>%ݕ�;Xw.� ��x��Ħ���T�����2�̓�?pm�b�:�w>��vSS����١�6�w'<�첊�#�"M��E%ؓt��9�����깈i�す������q�E&�N���C܍�8#��.G�].�N�Hb;`Q_aNj�[?��yZ��������Iu��a E�W�wK�v�kdL�F�a�t���3�,16��ۭFd��Һ|z.c�d,���"XX׍d�o��ä �{l5y:=�þ��n\r|�թ䟼Z�$�4r���n���H#��%,�.��P��������wJ��;[�͟w�w�,���n(
�$��ʹ}��Y�(�b�Eđ���ȍ�A�{�"i��r�L��s��+�GE	]�/�'ͪu��=�N�oyG��I>f��1���;��ɹmå�gzѨf����G��"��ӽ�Zz�W1ū+e�dKuY��k���'�����Zu� K ��u���ͭv�9�zݼV����KFW�7/�Z�X%�^^����y� Ko9�a���;oi�)��?����8�����H���)�׻�}k���������?8�|��*�m��2 ^0�d&`��=#�W|�!��j\��ğ(�_W�~�p�'̼����y��~f��cG��י��W�"�#�4�NB�*��NZ=>��)##���I��|e��c7Ap*�	G{k�\�i��&�~/q��9��.<׹�ζ�b]z|giq�yG�`2�;�_�t�HbO�_���� ��y��{o1�h%Bb"�C0���&Ȯ5�������}���M���le�����Z�C�^����K:�U���ܫ���Ѫ嬵���n��>�Cܑ�~�uT�^Cm�:��u�%�gLn���n�����F	%v��6�A�qEA�2���Z��������CA��/�4����W�����`g��^��I�Ű���C��e>i��%b���+�rQv(E���@x����~�����>O]�S~i�Z���-���35Z9b�}�a��Gb��SY��g�p��Ӱ-7�oW���s~������gkD�U ��j����_.����CȺ>�L�/�]���u�M	��H`�
��Q��|�Q�^9����:^�Ð'CL �W��e�5�h(��qz���L���sW+Z��u>����F�o�E����ת�3�`;�I:���a��Nm�C_�F��#ݺ0��T�V���eq���j���~��TX���X�P�:��{��"�T�54�DӍZ�"dYa�Ѫ��ǆBC�����׳x�3	Ww����l�@p���PǥMp++���D�QӜ����l�ߙ��ux��4x ��e׺��@��I�<�����=�F�����\���5r�|	����������.w����ǳi���N�93w���?�U�Ꚑ��ZR~D�:�L�����iK��v.o����Hͅ��$�ι��T��3!�7�7����sj��_�յ.�^W�@<� �Z��� ČJoy2���%TO��]�"���]��7x��o�C�؜�\���̔V�X���.��VS�˳��f���F�Sr|��:J���$KyG��3,@/�'������x��o
rgLI�������Ң^[[���������47���R�� '����;Y�`1-���$�t'��k׃��&9j�u��L�w�9 �6�nKá������� ��5�f���x>i{(Lz�]Z�����"��Q�c0�a�������ʨ|�Yk��me mm%5Ti���������!��d@�,���0��j�p�.�����G�:�?BC�*��~Gy�.�Ԩ�;p ǎS���ow|�Mիq�̙�fK��*��v���O���h{�,��.��fr�}�3W�>L��ė�52�vj����0�ϛ�����w2i�~\��3��Z�Dm���p��ȋ�+~zʜ�	ܜ����2k���9sRI-�k�����b>ztl7Vvʵ�
��;�X&@Κ��=Њ�f)�ܲ ���:}䌏�(�-:��G�Y��Xh՗�p����Ue��g'��9�ߨ��f�k�_���B=�[��V!B�duy�4�v
~qBA��N��:IΜ\���ǘ^s�����'��*������ų�>`���2OW�7ⳬ��w�� \���o�3@7��n��U���������!,�_@OU�-��7�t�>*�8z��q\�r�?"�a��JU]��w55#��.dD��x�D�Z�L�#�k���A�M����c��$L[4oW�j�1���H�4���s:c��!V��K��)���g;��{B4�6���cZ�A����n],;�vh-+ur����a�x�!�,3�Z(񁊫,��cz�U٪��^~�o
d1�QE_?��+$rM�adŗߗ�������8��.C��4�^������g|�2(�"��ө~�o%;����z��5���і��FP�T�E��k�Q�C�>��q��E�\f�;ES�KM1�3�����J��f���9oզ=���7������T��Է�xh�,�*!Uh6�"�>��ˮן �b���/�Πdǹ�������!��g���������Z"�:Y^����gei{h�m�����v��kf��f}yM��@����7�i�1���ʮ���wI�rn�~�o�lm�a$e����?
�~4S}��!���D��L�x��������;��pL���Cu
��áT o��IEA��o7��♀5�����޶�
�83,z�=�>�ap:�i�(��$�u��G��"��y�7��L{�`�=�Ok{s��������o�H����2�S'��IiM�-7��2��O��T��e����}8(�h��W2V#���`��
��e �kmR��E��G8�;�當v�p����D-�7����7\j�b��;)�$l������d��O�"O4L��g��X~A6��4��ĺx5�^��������f��, ��/�*�t�#�:̅6t�3���x����O9L&��^�!&�!���wV@yů|�L��,W߾�;;��*�w����cYnkJ��*N!�4!!���>!���e �M�ؿ�$dWhzֶ�� �~Vb\����n ���(�|j+\~=����&��O�ȷ%��&J0
��/d��7Z�R�r\�&� �IW���W_��r�J%+�%$��d��p�M�����h��� F|���Gџ!a�{�[��8B��{TE=�A� ^@J��H$efe�\��J,O��TspZ�>��\c�Sdn6/^/�F����4�o{$V�Ԧ�2gkV�>�.*�= �`l#�*C�ن�ͣ�~�	��]!�L돐�������3��y��m�܅��Y�4b��8p�;�p��^�hn������s�N����пˢ>}�};����}uA,---8���T�4��?�_����� ��� [�5\���5t�Wq����2��G��?����8�s�SMp�Ђ��Wq�?�B�|[|Ipp�o_�7k���L�V"];��I8h�H��(!�d��������x�BI���YK$+������F���ИڑJHH���jc	b1�Zb��Yq�Z�)�h:���G��}��Ov;�������LRPﭫ}z#��!.�ӳh���*��T��!�[Y�馜T}4;m���vsnhF�r�" E��d�IE��7�K�^��%�=��8e𹳡

���%�r���=�OMM�KH�`}���3���QsSP��i/�:��n�ՙ��#�EL������ �����\L��E����w��_b[�6���Ю�[,�x+Е����c937g�p��n�`2���qrԠ�K�Б~W�����������w�Q�	���ɂ���|	3���D ��z��3�J�^������]9�F�f��l�M�����X�_�ƽrb�N�J5.�P�9@u&��eGG�4UA.ۇ���tl��_A:_m}|���  �F���{ZZ7^�I�BG�.��o�*��Vu(p����ύ�V@��Y� PĎ?jL�A'��g��ot�Ju�'[��waᖢ�o���+(���I�+^� ?�祅�}��7��I��= ��y�t\�ߎw^��">�U"�x5!����j'�5�*A��T�͏&��_�J�������S|�<�3���f�X*2�C|��$%�ff����mU���ܠ���N9qqqvNί��E8�ܡ���
���l��&~!a~O3�7N��+rGCp(�e+��{��2?vZ����+�Y0�����V[m\��<08(t�������֚�4�ͅ���R����W&�|�U�a˷�h��E�~�Rtż��D�L�h�7�Rq�Q߼^�W!������e&��9 �+�-�U���/�L_S_���[ �NM�x�u���7]y��#�/����"��%�=&!�����7�:;��d�㣔FxUd����8q"��oN��z���+w �d)8���'~|~!�U>==���Y�a�RIv�@���[��'~����Y��أ�s��_���#�U!D�0|�c3��W9	�w-M%e���%��Wo����gRy�ܱ�UQV6���r���������(lM����j�e@Br!�S�c��pڵV���SB���8��W��U�O>!���C�X�C���ɺ�������X�-�2i2�|L˚���,nF�r�@�}lc��ae�*1�t�ⴖV�[k�w!�����4=�=���D��|�F��t�cDE2P��k����|㯞�ť=���2=s��7xG�,T�.d�` ��RC#!T/U��C?=��������ݸ�;]�B|6.�ua��G�1%�!��.��<��"3�^1țW��Jݠ��=ɖ��!��B�?g�������e (Va���o[��E遀X�7T�ɬo����{௣��`)'� �,x�:y���ʅ�iK}p��nR�,�~L�ǯiQ���xR��8����g��	{��������OM)���@�~b��=���,|������Mj5�@`J`���|-ZYY���������'M���m��^C��ϟ?},f:� �x@�A��юy�����3����=�K�.����Q���c��;U�Óc�{�GY�T���7�e��� �����f�^M���\y������Z�_Y��p�t�����Z��y��э�"oI���l����pN�p�_|���X�YGA�$8<ܥ��y����X�?|�`��vv�I��k恐�-�˗��[��_`Z���[�e����&�Gȣ,w�R����[]�]�8|����s��� �/>���,pN��ΰ5��"�����O~����W���ȕ�n������|B.8�.t�^2��}u�SVH����I><�!���qf���|��Y��B�qK|�k�cOoo�3��\��������=���A�����=�_be��	�T�\�K�.D js�ܹ�������g�ʟz$���=�q�6Y�yB?���f���r)�J�IV
L��	�����;	_wl(�γF���<3�<�٬>����S�&�4WX�:O˸)iM	��{��R�-�m�o}U�k~R��Ç�	��v:G��6��1Ǝ���$���d�7b�W����fɖ�l���-ڲ#��Å*c팷m��aL�J7�;&��%�%���o
��Y%�4Mݲ��54�����4,֫n*b��'������
:FV�Łu�T��u���>���7�����FNT�4]2�F63ɀ�.��_|B�
=v���3�]\ܧ�3�<��=oL����q��jeR�^a�Ƕ�$�g��˳h�(c��ݛ[�y.R�7�_*d(����1x��\���bLE��bi���y��[�sIڋo����)U�{\��<�D�f�E�����%V�0&q��e���1_�l�s]܄+����F�U|���8m��0�5["��C��Y�=ƷٔvcG1 9���m�X?�U	b�4WB��޻B�E��'ZO^��@֕t9N��7�@�)X&�X���%c&��k��lS�BG�n
�{'�!�����g����ʘ(�v����﬷���h���,�LUl
�jW����>�3�т�0ۮbӧ�C]�%����^������"����G�1�$j��m�%F���k�J�g�޼�y��OW����EW�F^u��A����nҥ��'�q�/,�H	��e�Sh����A���b\�w� ��=	�D)`���$��
�*n�v�}�����0�R���.���^]\��X�`���B��j��$�[wC(�rE0�f�I"���[M)��ö��f�u�M�詒�n�Y���������$�������Q�qb�/~�9X��iwн��Xe�d%$����?5���d�лŹ��i�2�����a+*�0�Ɉ}��������m�0N!Cc��Mх6������6
J�R�������'N|�D�I*__O���m��1��R�z�;z�J6?`��b�v�*M��EMlQ�l�Lٍ���8v���صIٙ[�X?c����@�p��Q�oD�����,�(��-#�;�'	�4��|�g�Ž����8n�/>�~W���o�h��p�j�ߔŪ|WC(%�HBg��Ԍ��tY�v����5�4ֈ�13oI��d$�`5����𲴻�������/-w_C|�s��"#O�9����9ޜ2�9�q���]��u ;躳�ŝ���Nt�- l���#~�V�ze�Z�40�`�>�ⴚZH���p�m���l�)����i4�#|�k����p�!��o��g��1a��D �9hy�eңS�.nv��wo�U��[�*��{����˷��W�$��a}�K�{��D�4DM�}���e��hl�oxb�iN#�9۷�q�J���+�ן�&�
x�q���l�<W�*݃$�~���}����hP��`>P�3��G	��B����L�Q�!�𺬗�_X�t�6�(�����~�;ɒn#,����o��8��K3;�������Klo8�?�������g*[�{zz��[���!J��,Y�oWO(b�a��TPEM��<�
�\[f�)ߎ��̀�����eZubE���/~H������#�z���0��5D�����x�@,�����U�w.��F�Kg�[�V����{�W��.T�]ρ�M�c33���Lμ�0[F�Դ�?��������i�VY=
A�Kr��}��ΰ�ta/F�~S��!=�:��bz�8+⤹c���d��C����p�3�M\o]��6��K�U�l-~�$P&Bˣ��/��Sɰ4d�nڢ��X�"�av�ɥ�DDZ}������o��p�_#�"���z��J�f����Rȋ�g�/�6��*i�T�/Z������?N�;�JL@J�c[��՗�;=��׎�@�v+����X���=nM�	��[/��\eRi�����s��ɐv��R���'�?k������X	�(�����='�z�[�@h8��e�ޫ�k������{��H J�Z���`�$�g����vR��Y�I�{�R&�\~�F[ 'Ġ��_�ب"ek�f��Q����Ge>����3�kp7�ƣ�����-�5�
5�2��}�\.��sED����|���?fg��F�Zi�+;�.JVD����6jn�<(!!Q�_Z�CPr�)�._���y��/,HE|��%E��8S����nU�8��yٛ��;GJ%b�R�4�c.�9���҇W?~̪���Ћ�jl]�p4�G��Zɛl�I�,@�5�`�Evn|��`QG�Cy�Sd��l)�&;�h�����c�<j��`ܧИB�����."R�>��i�o}�}`�h%it�q�e5ʤ)U�is�m�\]P����?�'๫b��5u&�����qǹȜn��o���B�SA���~��hp���V�]0�h2�~�I����g|s�sgQ�@C��P�s�݄�MFXtǝ|7�mm������:P4*�=�}I�2�~��+��$�v}�};��1"��Z������߿������n�������lu���P�ᐳ�{��=�����͝�%-d)�i�T���@b'W���BġutR���D�p H�Ӏ����S���!��[���R<|N�o���y���_�h��:�j�,��A}H�F�4X�����S�N&���k�eG���θ�O��� �-�g*n�����W��%�1l���c及G��ܞ`bٺ��Qz������<v�vke�4	���Fe_�ag�g��e`�q�>4�K{($}�J7����p&����۴�Ý�:�NՋ��M��0�ݧɡ�`z`����Yg{���-��޵�~�.��Y?��ez�7�<�+ڡ�(���T�iݙb��&'�E©���b�U|���������qN���wK���9O��U/H0lv��uᩇu��(�a�>���mnZ��)�
��iQ�'U�`�Ⱦ�%6 �Ң��"L�_&J�KN|���0�)�@�nv���76�g�~���������T��귄3K���v3m ����'t���C�$*����3����jt��x��E��/j�喐H�;����;fs+��.ƈH��O�.p|��d)X��&��1l0�-��􏉔�˟���a?�h�ne6X}d̟{@��8�O���dG�''��%	�(b���M���?�w�vQW�.r����B߭�o�_愗�m�~/t���O�r��
Q �	�x�0�l�~���E�}
B�(�ݷB=ل���a���>!
�C!���u�zD3ږ7,�#�Ӱ�ձ�`�4���Ϧ��������[���ĸ�B��R h��=FZ�����8͍����������uǚ!*FF,*��+ZN����\_��G=ǿx�&��a����6�sq)�D��8V��Ȑe�0?����=�y&����-j�o����>q^����̀�Y���h���}��9������#�ϋ�&=$�*����Qv��3�zw�� ~��>c|�O�ˀ�d�:79+������k���ޫ,�[�뻣dר��@�s�b�o���ې��A%��ג�V>`�0t���eo��:Մ���v_��R �R$�F�_�;2��Gv�`jN�Wz�o�yVu��>��@K����#��n�Ƙ4���/�ijj�����|�ݛc�l��|hI�pL_�+��*0e�RDYKzm��&�us�����-���.�WK+Us?$�dt�T  �;���~�;��2�}����M�54>�TC?��%nk�择�s[3�&�֝$���5 'W]gz���0�SA�J������8�޻�><$2d _��I������+zb�Xch���Z��\V� ��)hG�t���������p�y�ֺO9\��F�{
����&�[P���#`���lC�Z[�m���O9����0d��κ��>ql�H��ah�6���/Ҩ��Ď��֍-jDY��;�]YP����ǚ�s�h%ݏ��1S�AU��d	[�Z��7)�t�	J�vO��4t���$�����������!`���霠� ���B�}`܎�7#@x�#�8������G��7['��l��mؤ���[�"Y����w����ڄ:��}�$�[^;{FHOþגQF+�$���ʎY����ӱ7����5]/}4N���� ��L��d�5pfB�l�߹�3�ZW����PwR���$�W������_������d"C)��#~�\V�|��&3��
~�TvHy٘z�v Z{��Q=���o�	�\��L}N���7�|��87'�Y�����m(f���o��̌��.u9�s��x�	=(%e���Ӓش��XN���a�؊�@F�%,��X�~'|�A$nG�OE���������_���:��=c�j�1�a�8#�S��b�]�
6`��͠-��<_�[d�@�p�I¡@,�y�x��l#��! ���h��W�y�x��q�� ���g&Zc����-(f���K��%�E�(���
���> �_]�5 �j�����6!/Y)��  �˦ԥ�zߠ�-��s���0��s��F�A��]�	����2�9���(<2$�����$�>���#�N9�ܡf�7P|ے^ʬ��t�9DX�o�l�V�a��Y!z;��{d��,��	���<�&�a�,����G�̌�F;�f+�|������W޲��#G��]���£+i��0��mk.������؏�
�w,�Qc2�%Nb�TY�u��xvq�"�-���O`�;N9�$Z2�M��� �PT�x�plZd��U�A��^��@�e��Sy�>�\|4��Z���]������Z��p��¼�%H�k��#�K�#���2���A�;kc���8q"V��Y�Ȥ+ �T@N(`���D�KK��K�
a�<Z�)𒁙z �>ȅ�l�A��
ԋW�O�:?�Q�;k���"X8��7�T��{o�WJ�t�Z\�;Λ��M��ZK3f�ִ���3��if�G�/^��Bzl�U��ev-� ?����p2B!�i�4)큍��_�&!CX�z���o��Gggg�k6?2_~x�lE�#a讫�����Jڥ!����x�Z�(Z��9��g�ːF\�^�N_��߽�ʯ��C4�X�z��F03��\�������*������h/��I�)}S~�uT\��O��D��J��>����Ȑ�n�\�9�X\Z"]��Y�휀	 �A�%���܂���1�+s����
(�E*CP�#*��8b|$���)�`g��<��mpʀy�(�-4׵k��+��k��.L���R1�,�;��ΌV8�4 �ꌋ�n�� ���I=��~c�'�Pw�Cg5��u�6���"�<;1��_ �u����+�ƈϹ�{`���\�!����}%�\|v�ZON� ��4�����%�R���
v��Í��}^^^`EJ,�
E]�x4_���P���
+/u�<�5x���'n�P��A�s�5�X<6�N��Xj���ܥ �t��I���Z��2��}�9>�߱9��B���ZfA�0���M Yg�����㻙C�AM�O����0ֻ!3Q��Y����N���*S�����S�崲Ut�.���xY�]d�h��53�:!>�T�a�ܞe3����0�%�Y���k����m��k��c��ʁ��в-�"��-q�4oP�<{Y��$B-IL�i�o����n��B#�Q{��w�w��6Q̨���:Cat�J��f%W��
}��Cx3=|����V��|(��t�:}\ՙ�0���o�_�fHI�}�n�y�����~�*�:������V��雗���sr;%ԠU�'Ӵ�ݿ�H���g\{lrz�<��rD�W��ݮ�=[sL�l(�?� �.0>>��ɡZ�|=��!��1
`�֗��)J���h���}�	���L�6�jeic���A)w�Β�4�¦���p1x��ՙ��R&|�%,�c-;�����M%���6���#l��t6u�lC���ek��ѨZF������:tsI���
��g!�s��`���3/䗆
�r�wtw�H��`~�(蚾𜘜�E���dw�JI��Ɇ ���`��S�K��21$��"�+�+s�l�L�1�"���7ϐw��<3�|�PS��I��38�����δ�6�w�E������]IV\x�`�dmQ!�1�n���X�N������x��x���ϊ&�CI��Pz~�A�ON�͇	RE8�&���Z�o菞�څ�ʩ���ve�/n�OAW�WԘ���j|wo�ﴥSN���MK>�>���ou���G�WdN^��`a�N�Ğ�b�D�l\��b䃨���]���Q$����˻eu����콒��b��U���4�$�I�bUt��?p���_��,V���Ջ��6��1���.jhb�¹�������g�+��Q|z�D#8�G�n��}F�����_�\� �HI
�x%���'s�~��a%�
�FW�N�U� .(v� �$�yxZQ�=ub�£}�q���%���b���d��E6ZZ�ܘb��keӛ�ng��,,(wt54hzdJ�7&���E��w`�8u�C� �h���מ�� �����uz�l��c8�@˓G�8���Ӕ��8�"��oq�<�9-�v��$J&���F��k�U��|��������v$�vE�HR�,�![~��R�;:\�zj��v�a��ާ�
GA���	8B��W�ѣ�V��L��8w��y!���8��%\A͎r3�>f���{|^4�L�" ���w��/`	����|��U?��Fœ(X�l�F�/�q��z�q������'����K��v�!U�/���Lv��)�^#����_��X��� O:�F���uT��@|�� @����S�D[�h��Zo�Ǳ�J5��6~а��Q���= �`]�N�����.���y�䊸���u�kO�'w*��g�ߦL��O24Ԯ"��ԣȁM�Y� (`�_����h�!3��c��=���'�D.�zSa�b�7���Y�l�2.�_9I� ��I��g��(wo_�o+z��2hR��ө�U$f��@��Ǫ�\ǜ�^�V��}��f��]oAu�O���$�73@ɰi������4c�5�D0�`֛�>�8���`WUU�e=�] ~t?s|J�\�q?���D�������f9��1#C������|�����	Hq����i����U*�����Qsx �[���':m�Y�����D��1�,ug�q�K�����6��F��Z��y�/����n'� ww�b�l��6����[ �QFO.�#�M��w*�	�q#S���F(�v,���X~�U��6cĆ[y�v����9k�q�h�ڱ	�)_�2^{Ӝ��vŨ���Sm�̌Y�9 �Tj������؆际ezI���_�����A@1錘~��/��Y�2Fg��וme���|1Ԗtܹ8�+���~p���Ҧ";_x�T���Ė��R������*�W�&���PCOI]�.iH=����п� �V�Vi ����o�-ӹ�X~:����J�(@|	"� F�j��D�Yn��AD.@�}6��;��Sv$��0�@�IݧM}��f�~���ie�ˉ��v�ӯ6S	*B����6��3bQ>>;��/Yo��טlQuwO4־��-�-O��݂���<����~Qfwɩ�lB ]6�W��%�}��<$�4V�_o��o�{��i婹�V��D�:_�Qu�Tݤ:j B�+EΦ�����W��LA.>�$����v��8�r���0���ߵ8D��@R�}r���g.�~~��#����tu��7'�E��ͲHIq
����>.+�Pa�Qq���ގb��b�8�cd�co� A�#lc���ґ��Ȯ��r�T�1��{O�ಢgZ��*2d�F���ֹD����4��a(�,ҋb�K�5��R�v��=�w���|v�&�e��aG�O�1���s`�����������	���d6�W��4���:f\4SWY�.��E�5]n�]Pߵv,%� ʨ[c�kWQ%�9 ����l4�rbf��1�bڼ�A,[�FuTτ�.��,ԙ^����� .>��lg�dB^G�V";#G=�J��	 ���aLZ�Z#f��W���T�o2�����0���TN���n
ylY~t���0��4��'�[f����֥cOE��(���OCCn��,sM�R�y���	�V����h���0�	�T����Ûw||j'�Ͷe�D ���O��O������N}�oRR�$��~�;�1�>�>���r�~�����L�WW>�y8l»G���%%�J���!&��+8~����	�+W�(qϾ6+S#r<vWW0/np5�n� e��_�b[&�	��#��=c��N��'w!�4f������`�H�@��kh%H��Ga��}9t.彻сT�V�˷���n����t�9�cv/�S��i�	z- /�F"�9��j�R�]�T�_ff�B���?	�£m,Oa.))�GO9�-p��_kQ�Q���}ؓ�AI��f[p��%�7�K�P�z֥ގ����b��8B����=���'�~p�y�B�}f ��e�S�-ش%e���.�|���cM]�æq�KZ(����\���}7�Ě��2�� z����S �]�GFV*��h t>�=��e�gI�<�k��?#�oΡc����}�6�F4�w�L"� �'�5�(N���Z��Y���Ŝ��� ���<R�<�M����yh��ո>�,�����ct�:��w�����ߞ�����e��q��SQ����k�Ӽ#u4Y/�����C��!�&w��˜�wV~H>n݈sk'Dt�n�a��3���1Ş���;5�%��q�ysl[Nc+V�T
�j@GO��"�	p����$���x����q��8��Jp�,K48��}��]��c�c���(�T;�Zذ�cHܥ�f�ۈ���	;�Ɉ�6�v��g~d����]0ŏ��TP�+�i��<�J���`���9UTT)n����ނx��l��tދ�BZ��^�_wˍ�Ƙ�i\�5���X�j��q�/���4�������և�����e�%%wq�b�*c ���x���=Gm�Ej��я�˺�lj����T9�k�R�"��~��A/���K�¶eV&^%���L�vbQt��l�d���KD�kՇ�fF��w�a�����TA�T蚵=�|_Z����y�{� &���/?l�օ5����F����x	BB�cIp���1�A��Qm��ؿv����y����5�NQ}�W�7�؄o���O��qp���j�<���4�hJV�����_�?�:�/�@�;�m;��x��gTN�6b����HJ�L5�y��$��bk��������=淎��K���z�ؿ���~S��rׂz��/�Mk��Y���_]��nZke��@�Uo�?�V����ҵ���8cV�l:O8}ʉ36l) �tY�Wf�^��Ԫ��Ӭ�FP��x�ۍd�|ч��t�/Ӧ�0�ٷɰ�ҁ�ݲ�/��j���?���|��R�h��;����7��m����'�'���a��|Xp�;��2�^�D�br����W��'0_�L�Ԭ-4�߳ƏE�n��r�:��xO)l�Ma�6TsHw�ڢ�ق�Pt�j��p�5D�/�k��ˣ��)j��_M�c;D�&�G?��,�Wۨ�H̞#�r7���$�r�Et%˛w"G޾|�RUm+  �(�ƀH��X����e�#�i�/���aa�0I�$��,ǋ�sJrӦ$!�y���g�N?$m���U�lE���꫊�;�s�J����d%��䍶��Y�w.��Ά�l��m��#�M�t�<h$i?-^���G�JSl��/\K;�!aZ-��aG7�;0¾��2oN~���z^ �GJ��ޗ�<7�vj�Ν��
�9�Mڋ��M�F,��&�����4z�E���*��������]%H��|��Q}D�I�[���Cn-Ն&�4ern-���v�Cu>*��3��g�.m��:34{/+o��yv�k����xh#pp��8p`�ZGO�W'{v<ʰ�?�����v�pIR�r�d���ˎ��U���y���9��dCN��LB:EI�z/]H0^����V�,��O���n�F���x��G!%`(��:6���aL��L��K��`��s@k����zo���щ���ׅ5��	�9}d)/�fG^�{'�39+�+x<Y}bp�mU55��.Vf}��Pf=E�0�G"���N�>��x����:;G�^q���Ge[���fB��m�K�ZG>d��w��?yd���L��/y4��ϟ*�:�>!�SOYީy�K��	����� 6I�z�Kxm��נO�90䥔u�|�/�]�AH��(?ݧ���U~_K�P��+Z��mK7�L'ߞs٨g��C*�'�+	�n�<��#�>hPx�l�|І�W�_"��ذ^��4�����un��O��宾����x�˗ٮŹS�ʩ��Q&ݩ�n�g�3����~���A-���Pߛ!qe��j�
b�ظ��!�n����7��w���`hY�@�g_]M�2b)Fv��}뙕]���:^���O���p�$�5� �F�����j�Nr<ʼ�36{�lGa{"��I�U��]��֋�՞9�~C���\��a����M�t-|��	�ƾ\m~�~UQ�?+���a�ѹ��I�>s<��NA�V1&�Y�hhe]���!��ϟ�dv&Y��%�]�E,�	��h��V��%p#������ l�2Q֞N�vfo�`��{x��᪤�<{[l������wd����ܘ
 ��#Z�"��	O2� G�>�o��,��n�v~�+���$&p���f�c���e�+\Vo,C��)r���X�ip�mo�/�wl�����ϑ��:�Ρe�`vp�J�Fo�a�û1�KjV�jv6�ua0�4}f"��Y�(~h74��8�{�	��YJ4��ҫܻ���*f�`���Sl+dQ� ��?�Vv�m_��D������G��S�cL5_�Q	��;h��2�j��yjBl�o� "I�@�T���׌�;u� )�VK�n�Ȉ�k5��+�C
�
a|f�ټ��M`p�ofR��Q�f�vr���X���A����_�A� qn@�������8��fb�x�;lXB�S�'�>&G�����I1�,[���_�!����(6�,��N���B]��ů7�g�c�j���vr�+������? p�9���GL{Wp�?���y�.SG�~tgn(��q-2n~K��-��B�ª4!a��>���� %��\]��u�]��b���5�M	p�4���뫀����j'�V��j���p����\�Oλ�w���$GL�Sy �B��K�{��>�2��s�h�:4��T����3��hEm4�����~�9�%^�y����b�.����*5�w��]��]���z-
 ��U~�I�z��.�r`A"q]jM=1���}��,�[��M�gY*��zQ����ռ����::Z�����Ʈ**'6�73q�1)�a"�ۈ�fT_@@��@I��ޭ^C�&F�gX Y��NыV��v�5)�i.�j=!���O�z���/�����4�j�3Cc}}閘���ϣ��k����؂�ǟBA����ď�L�?͎��1i�:��|p-��t��=�~)H��U�W��K=�'�t���%���y�R�������d��O}�E_�gr�F|>�����q�PMe��p�" h�i�ET@J@zD�(M�"�)R�Q%4
R�H��:��@�&�B��E�����׷V�JH�9g���]Ͼ��熓��G�;9kn�u��%U��V+M(mo�t��-�V^S)�;	�}����o*Av!�
��� ��!`��M������G5��N�a����C���=��ֵq@jn��DII7��Ve]ō̚{�8��r����J�l¨{ug����#���<2>�>�����x�1"��|J�5���`B?�=�>���3���^�U%ە��dz�G1��~�YOKnU tU��-��׬ͯO��?ؘ��z��e�{���TZ���'/�V;�f�]}{i�������\���:���/_��+Z���a�l�9߽�p9���܍�9փۏlՔ^*8�����7C����&���*=���c��B��\�����5��ɘ`W��翸yms��&o�?A�z����Ip�MݛZ0��(�+��f�Jk���u���[���n������'9��M�<�.����\;ē�(tF[��6��ԴE*)��%*�m��kY���y����{�:V�6�V�å��i�4�.Ch�W!Č�3�I:�Mn^�ǻ8J*_��*�)��o��g�=�����T�Bki!6��׼�0b� x��;$�zf�Փ*�7S4�_�IoxZ�o2`�*;p\GCb�t��h�}�j�5�b��̋���o�������g�6��/�(dm���m�]*��_.^yC�]�.�<Q��^?�2�-`� ��$�u��W������n�����g���ߗ΁�a>s�"��Q�!6PDPg`�^�
9G�yM1�"�!7O��P�1T��H��J0�Z?�"m$��z�3�bR�n���Z�?i\�vi��u���KNp;�N���8>��!{�`C�� m+���p���Ђ�U���d��p�#_�,D�r�Ƨ�oe���D/(9;�1om��0V/��3��/�����p�ݧ�f��3<��C���� syb�xT�e��d�
�
yf�E�_y|�Nb��CF�K1T[G^�ϛ����!�&kg��5�G����P����Pjv�L,�����<)�>�`(�h����C���+��x��8b�؋��D`�R�:#�z��1-�YaY�[��D��*�!*��J�S�	I�����!�m9� ���Ye���������_+Z0)�[蘃��V��L&�I�Q'�,|)�X#V��&%�r+��-�{��Өop�5ߏ)~HK��]��\�ih���?vg,ֆ�!o�����g����{�쐗wԭ�΄/���OM���#wj�G����bȾe�3L5M@V�IF�}:$@=r�N(O��
W�I]r!�,w)8����|���v")Ο8gk��S狙$�K�3�3�l�@�LOjZ�����%�^�h�&f���� �q���Ew��X�?�� �^�l~������~����G[q3ŷ�;����T�l�|r�y�}p� �
�`�f��zZ 2�M�m0S�籩�}T����DP�7�{������tZ�\��+�Km6�!TjM�`�s���Q�a:�$�jz��K�h|Iϙ�+���$z��$c�?�[�k�����ݻ3q�qk�ݡ�B����]@?~����p���������^m����d}Q��;[�;��1u8M̢�k���.�ढ़��LO>ë���?Q>K��BFl�\�RJcq�x� 1j�K{5��~*\��FT����ˉR�����75��2^�#I۵����*y�u�ȫ�s���Kc�Z�6����~ ��y�AT(�:�U�-(܂�n�#�� ���zw6Y�at�0��Ҋ�������Ƀ�JW7�	���6�r��k�y��>;�(c���֒R;�gv"���f;zB��r"��3�~���k�>�Ec��=Qx��*+@;�eφb��Mx?�q�U�t��ĕ��vqV�'JK�-N� ���H�����ّ���	[-��?Wݐ�s�H��h�9��B�8���FN"���<��W�)6���e�����]Ρ'��VG"]r-��zfanZ���3'��R���9e�A�p�K�F�x/`�eJ|Y{u���^��r��KiGs����l'��e4y��q�Æ�f��Z�V/zG\()QN�?��x@���k	���?{�d�6�`z���B8�G�ȡ� �$ٴ�1r!�]=P�s��LX��P���)�6�£m�?�6�+��2�֬޹C
�N���QpI~�Qi�'*�\ښ��)�02��YO���3�`�{���(g�o�N*ެ�$�K�Eh#$A+A�����4�%��ŋ������N��;���b	O���3NQ�^V%�U)זҠ��O�#hMg��5���T�u���N�ѱ��E>8����Y��|f4*��}����P{�ߥ�$���<��<3;{'��x��eDΩ73��ͯ[����sU.�G^n���}9qXڑL2���7���)]�|��+z�4p�Tsm���Lh�Uѵ��yy��� ��!T�nU�ey�౷=�M?���LĂv�B9/��h��nلo��T{SQ�?�n��eo\����cA�l���5�O{�F��(X�_	��y�%\�r��|�qT��w��T�1�i+v�xX>c�rf'S(z��ό���:\�l�M"N�l!�+�n�q]�%g��~��o\A��ǩX� 4��Ў�R���.w �^� �ٍf84��F#���,!W��t-�&��t^����*��mHL�C�w����$3C��r��yG�x-B������#�Ew��U:�T��gpi^@	�+?h��}�b"�t)WZ�N-�>��"�Ɂj���VaҎ����~�k���r��������G�o$;�8�r��*��tҳ�l\T.�t�q�_�q��bHc�<��K��d��4*�Tׇ������@5���r�,vk�Bb�@�W�[�G�Z�C��O��6z��� �	X�xP�{�!�?}&'���8g���8���`�j�c�LR=h�[���ʨ�j�B1jv�x�[�[G;4F%�Qʪ`:3��D|�b��XRTM���q�����J��/�#B�� ��>�K�cS-,0��z_uv\,}0�H�6�E���D�-��w�ޜ6#�w!�+4��4����6�
u+1���~�)��r��=� ����5ggni 1�|��sJ��f]�`1;�V�>�#� �hx���y������;�[��9�����������]�hk�a"t�R�m��v/3]o4�]�ʹ(�!��V��3�=�������*q���}���礐��r'f"6G����K{(��N�gA�2z��e4M{9>+��nk#��dP�R��x7P^��g��X_w�@>\[-��4��.
Fs]����Y�i
7%Ӌ��h��>����"��uo{'�����a�+���A��e�jX�Y_pr{��l�%�t@*�4}�̪a�t��K�~��EǲS���<���iw��x���+&#���
4�[^�8��B�.չ軝��=5�ǭ��BW�^8D?n�wSݶ�������VW�bՅha���]���x���cP�µR�B原mE6��>z3xS�^�%3��:�S�>��:�A�g �mL�ܟA�я�G������6��Ӧ�C��h;�?�����B]ѻτf�Ue��kX��h�F\Eb{�����^Ő�����%��Q����_ԩW�qI���,��v{UY���3�|��R�f\z*�UR
�"�{�I6c7��'�,N�mՐR���Ԑ����A+,ݐi��O�-�}9�P〩�+�;��zu��l��{p��h�@?�7��q[,x��!Z~J�~S����
s��8?��͎�t��ȯwt��v����}We�uL�v��3H|}� �9��3���7���1��r����А�� xɂ!}��]��=!RI�U�E~|35��E�}s^p�LY��в~��f��5���uE��ř����n���Z���v.��v[έ+ږ�/���D�{��ٟ�O6Psl)r.MR�|�}�Q�������-�&2�4�=��M�ϛUڄ��-��!��+_@��`c->wD�^,�KL3����=p[�t�?m9�s �H�ǮeV�J)�.�]�l [m$�J�N���_D��\��j�`2�4��'��.�`���|^�/.����|�b�A�`�'�B��w�ƌq7W�v @���O���ہ�n�QXL?��ϲ�UYYY���p �yw�9��O��Q����^U�� 11�������<����e}F}�cI��un��V�5�X��/�B�C��o9h�ֈ[�p4��++���tdY=��(����i�c"0�iA����>�r!�Oo����^��.#�c��H��E�A(�k_�D�A� �����7*} kaR�)�.�$�{�������/V�꣕��Y��c��ҼDZ�E�B)�a?|Xw���E]]]LN�]���}�)���b��M��ST{x�4;&�T�׎�џ�Kߎ�ݦ��Z)i�]Xӕ%�7ӕ"U�
��Iʝ��$�B���4�j�������US�g-�-�������_X�_h?\�Y�$X�H��;gx*ul@ʔ�6��ٷ�a���0 ��aR	� G���B��-��BfL��6�������^0���u�	�?�a��9?���9����-�!�\�S��!��5��!��O{�X伔У(�4�V!�Kbs�}����Y��)���Wx��ߗOn ���s������%l�>�KBSz#1�BF��9��~��H����e��d��l� �C�-1���hx�a�����]60���|w�q���l~>�F��_�Mn�P�������4'�\���cO��*Mf�C"d@$��3��E� �'L^��-�u��5��d2y�RO��X���o�T�@���5:����-�T��Q�2D94�d`����e��,w�62����vA�A�R^�/�� nE���Sq�i����m��,2j�~��d��\�
�63��u����:"7�������ʭ��䳲�E��Y�6�+�Xr�^�7�O�>״'�y"����tvC�>j�^���/��ᜪ��!�-5�O>��eY ���Sp~��~�{����u���OT���ֶ��X���-|A��Bq�_�3B�k�ٿ^~QT�[@M!|��
zz���2a�eX%0BUZ`LB-?��[YX���ބ�r���EB�8�����k6}���kw�q���v7�f��I* �5 ��L�;p�i#�J>�[��6���J;���_Ó,�#l(5ů̠6~�ş
�
r�&��2�%�S,��E��R
�|9ƘoYy �R+�,7~�5��þQ�}(a��I�1 y���x��hyl?�(jU#��� �\BJn�+^�P�T�*����~�I�L�6�El��G���	��c���:ƃ�Қ1������w�c޿�ɝ��|��mA8�a0�w��� *�+�4�y7�#��^�������w̒~�y����xNC~��7������3���:?C�b �2 �2����7jT��pP�F���\�{ 52 �{��fv*�vt[��	S7�\��D���M^x e,����X���u���4ސ�9�qW�� �Xs�! }�te�+\`g/�{�32.����h�BF��W����+^7w�7��Ҁ��d\����V�$`���m& ��A�b�"�u)g֭��z\��+��.!�y���Es�$�H�K�yu�Ŏy��p"�HⓁy��<�x�$b��/v��.�q�hR�v"��n�t�qT�H�[g�a���6�ZB'0S��Ư���!�xaސ&^�[�('�0;�+)m/��3���`�@�,��1 ����N�ǭ:��^4�	'H���'i��X��k��I�3̔Mj"�/�ȞA��x�ͩOB��G��'7j ��U�(�M��� q�^!`|M���4�Wp��|�Kf�lnmI-�}U�SY/F�9�����A	�$�[��^/�.D�B3�����_��hw�N��8w������nj��v��9�?�M���=��F���L�jC�>�εA��	�-+��S/�ݢ����^^s3�6���v`մ�(4c5�d�%3�?9�4�r���C�ӮC�.e-NKK��$�hXs d�y�ٜPƾW�~˨@�N�h��,�
yZT�}L�w��>��o�R�Y�9����/@��Sh�BlPW(�����L���2�^@����fdW��/�a��½q|>
b��I����I���'�a 0HS�����Ò��vN�gH���=�q�����A�܎k�Q�Mv+%��ꓓ������a�u|v�����g���k�����[EE�O�Sw���EF&V���� �o��")N����|V�����R	�{�A�6��G�����y'�-l`��na[x ��,��	�{��s�
�����&YX��:,q���#T-h�^�s}��̤�P��Ċ+�:+W�޿7(F�\���ΪQ*�awo�ƿԼ�����k˝|��+_L���3�F�8^Rf�(`�p|;�Y�u�J�!)I��plw%��g6���TTkov�(�#��~XmL�NJ�G��t�p��y��Mu5��C��K���N<�Kx�`�|�Y�����m�J�]`��p�+�m�jc	`��e+���S!\�)�F(�@A���f�6+��if�M�;s"�/y����\���g+?�n��������sDF��u��ĲY�?u�
���;"!qVܢ\�2x�����?�Q�3��؍��|��PYT�0�N��l���r��'ۼ�?�@���%d�v��ۈ�:��Ӛ����Mj3�gK�ڗ��-%�8����I47����\��<��7��#b����8��yc������P*:u���x�F~D�}��2�H�˺K���e��
.	��\��AS�d_A����"�A�����ɹ�t��m������"�R��>���7�����!~�@�.DN!������-<���g@|f��?��=��^�A���ց\�j��RA'-�@J�� �%C�q�k���E!z^=�A�{{�zN��S���* \!��)x��sE��k�G
hν�݇���V_���������c��@퀐Dxs:H�c�N>|�eB�нp�e�rrG��$�\�v�^���ѓ�w��5`f4��!"7���?̸�#�������1
K,��6���'�_JژȨ������08(l��aˠ��!��G2 Mŝ=�=O���7�;�f׻��6*׳��W���5������l(f6����up�Q�e,I�q��9��҈h��]��}�4n�A��R��G��BmRY���� �[-�C�#�%W�M{օ���=M����Ƕ������:�dg��\�i�؞\ޮ#��������u��׋�n�3n�_�?5�:�ަ���6�h�����yno�x���jeUU]
���P�A�3��'�<�&m�
�I�hrOnm,3G�T���rMq����� ���3�<�� ��۬��᷵X���9��t���K��~�7�����T��sss�N�&�O�wz���޿�W`��r�E�Ţ#��*��P�%���T#S�<NcK$�'@�e���� �����̥U!��[[	ݔ?�z�pR�d~��+_�(D�͹Xa?�9���B�����#� g�Y�b�#�(��y"�E�e��^gQ�F�E�����߈$\4H=����su	��*�أ=w��py�Vm�k�{�0(�9]MM��^E���5��q6@�s���N�%Ҝd�4!c�;��)����"q�jr8�HH<VX�L���8M,+�u?'�0�;�aP�����qpPq$l���8Vˑ�5�Эi��5��|�AMI�(���2� �& iv 5{��7�t)X���y�_��6��if�>�����Yg C��Վ��R��?�:�
.�Oy��q�(��U��R�S�
�C�l��&��^y�ÿ��D7G듅~1\G�����1�RK����4��1��磼晄�j%BJ�H�+u����=���3�C��0�����������_��p�	��KI/�ݩ�1�ޘ��+_�����V�pTa*�w�6�)��7�y/ou#J��!��mK���F�PA���j�AJ,H���l7wZdS�Y�B�%
��^D @dQqn�p�����jP��e]w�Ӭ~����dr�L<)$��Q�O+t�ԇ>y�����M���&��� �ޝ���7>&��
&�����Pl-�������H���Z�͓m]w])�`��A��T9��)�U� VAk�mf��~@0I; wg�Ơ,��2.A��y��	��4υRh��J��H�V��lӭ���ʷ��'�B��F�d4�wIjE$)H �jh�z����	F^r�^�'�Դ��4vp��F�EE��y�\0��G��y	�X��8z��W��[��P�� �)�`�D,�z!خdx
�7�p��a�
|3���D�; �҇��H-$
�JWX?a���Y�sT�W�e�(�R�ʛ�4׮$q	#�q�����gH��\�~o�qP���y��P�)�K���5�P�p�)1+u?�4Uj�t��\���UaY3�^��q4�W�N�wjkw�=�r�<.h��(l���|��F��;k��b�'~�"S������e.��@z]bS$����G>����.Iqs:�)
-UG8#nS1`��k:�sE7��6�?���W.�
)J�[��4�E��?')�ut���[)����>,����&�i툼���y�+Da��HR��b���+ ��쒹\f6:��1d�6dF����0]�_
K=y�G������l�����>��o���&���B�C�3J��J���\�V ��s\w˪����C���:3Ǒ\CS�Dl�A'���۠�
{��x��0�X:\I�3J�"鴲���r�K񏂆�@���q]=���ӳ�����0j\�+�bN8�"��ʤC�+hc�q����H�D�Ir��;z�?hDm&��7?�"!Y��^%P��}��f/k.q���7^�r�jw1�7�����ZSAvI�ˡ���u_������BQ0�bx��MNb4,�Aԛ�X�%a軃睻��p�9q�n��	�<���1�i����k�9��S;=��	������5U]-�����&��^�� �t����'t�c΍]å��'e���Z�>?�pl�u��t�V�.�G�ܞ��O����|U,V����$s)q��Wj\_���pV���dڬ�^�`�+�n~XH��? �ܾq�ެ�B�`_w��!ו_B�0�t�����
��)���Q��!k�����vK�h���_�R�Jb���>��ʵ�[�u��\݇�l��^��C���4I���n���7iQ�����������0H�J�����l��-0&��<����BM~�$/ e_��U��b:RٔT��Zn�k���5��/]ztTR�}��,=�q��o��m���	��=y�ߓ�ݏc�	+�L^���3oݺ�F��^����3L���A��X�(K��� ?����:YA��i��5�ߌDZ�^@��Y� �+�
���eo�|0���@��n�����u%���_��_���[�3��JX��M�Ł%�7��d4�,���hޑ%��h�����8�e�C(������tN��e��Ug��W`d=h~�?6�ԈJ2��!��a�&���g�k-`e9V�r�5_?��j�}�2�`����4��D�/掏8���%��93��m�@��R'�����6?`��_,+o�q�+W2�K�-��{�Z]�CE�s��d�4ʹ[e5�&bDG ��M�mw��/�>ǀA�Nɨ��	,L���������.H�{�_9p�i�j�ہ�$�(o�x�᧡�3�k����%�
ֻV�ü�w���rT��)(R_�; ��jAl	��g��N�a��������,���Mzep&q*�����ޗ��Ɂ�ot|�����6ߛ���]^�ԙ$ф�������@U^f�0-r%��B�#<xP�=T�*�C`�\���2ʊ�9�1�������mf8�Z���K��i��������	�����{[Mj�hV��3�(fe�����1��7��5o ��bWݗB������e��&_{��������`��<���$�W*KK����#�r����N6??7f��X�IkȐ��;~s��l����,�����O댎��`����P�	i:��x���-���O�=z�i������h����
�
�ɜ'�'�Å���ǻ��d&,���.���Y�q���Y�ה� �H���FC�r���]}%.�K`dO�ԩ��Oi�{��p߱B��=���	����s2��V�`�/���:�g4G��礝(�vHd�y�*�q�Ю
^�v�����)M')��7ov�d
�	�nH��g�l8t �N?$O� ���'�E%.#��s��� �}1 ���z�o�9��C/�"�����Z�k����\N��|�,,26�$l�<Q���;,�!��Q�KƦ����0��h�h2p �AQ_!߽{�o;�O*��zg�ц#`�B���r/��9��z�t�WES�ޢO�����C���c��PkđB��Q����k���"��44�k�7N�����R��Zj���,��H��9�J.^I�\]��e�?�5������{�m��·�$Rx�b�s"�.�x�a�׮q1��5�~+��lR�*7�9�Pp�F�=N#��e�6�~`S���4|,�%����*3k0D�KE�d^��V_YXX�h���dY���RSS�aHW�Bh+K��y����@!E�'6��]iJ8~�6�haO�y�{�eεht~zPܣ��8.�r��_`�yKN/� �ٜ�./��:\j�E�}Y4��k-�[�$Eû� Kw�c��K�X<��T;��)`�fP{����-11���a����n�_.�	����w8N+w/D�;.f��׾t�7�㘟�o�t�7�>�z�oj-���`�˃�,gϞmX�D)�u��x���1�Q4��1�idcχ�1~eE��,1$��_����JC�)_����d	]g�)Tn�(#|��} ~��E�ő2۟Vg)����ô�\�(^_��p�)�Ժ��|X�hSt=¼ġ��|cu��U?vyF�p��]���#bbb�m����7�Ǽ��b"a)��5�m��l��]��u..H��)_����yƖ�v����nMvc��-�Nq[���d�ޣ-;-������L��bb��ZO�iL<����`���c5�7�O�W"��'�.���96?s����hx�[4;���m>� o�����L$�[�?='�4v}��"�,?]�G�9(&�"�]���uW��T�XA9����}�f˧_��\����<���M�x���k��\����d�ג0;���Ib\�*���ݜ�C(�o4�,����[���,�[� �Q���|P�{����z���v�<`ӛ�H^�m�5;���~5ntD�ݝ�:�QY�=�	�
x�\y��@��D+�u��T�@?�ԞX�t��\���>+!�5Hw�*ފ~�$F6������>���Lv��>�������͇�{�H$��]��S*�Jv�m���������2DS���dM�z�{�8���5�){P
�?=x!2�.��1��7T{��+�w��qʐ��7�-w-�N�p�@dS��^�
\7�7d�U���,�ί�	L��m.<Qr�A^�Se�A��k�����8��{,�U�h����#N�g#�Et�S��2����Z�-�;��H
T+xى�Fzn�h�l�&�U��f���ac�y�+#UR폸1Y�U���WU�%^�W��+s�/9�9�/ޘTc2�|�Q���Ψl����?b��Ț%�6v��蒨Qa�̰S$��W�{G�n���l�)��5���5R���v��z6tK	�g>���h�P"0���-�}ٍ���Ak{������A+���>����Q����M��-�_O�Ꮜ�4� _/�z��T��޴���OC�d��{{Tȟ/i�M(�0m]����H#?�[�M�ʕ+�x�Acdn�G�vt��}�5�)2�1;뚧�,�U�*�H��2�(����g�RǊ��!=��;{�Z�`�>��4Bq��V��� �����jx.�0r��ԛ�"!סpӇ�R!��lJ�rW@�� �ݴ
�la�je�0�xtR,ˢv&��+��`��q�F��n�b[7%�[��w�����?t��h)~ut��4�$��_,��+D�K�;�>�Qe�5r���{G�I�-�'�D`���"����/���B����C��~s�4TL�-��o��ۏm�aS�����l�E=:��-��'o
�"���[89�aZ0��u�Ɓ��2�|�a�ϾRȀ���C4&Yٹ�$$������:���(���M7���9��ʯִa>�������O�d
�����rKm�S~{����>�?$t�!B�C��6���+��ՙ��:��WlZ�_�������9j�M:�(H|ޕP`r^yS��/�n�� �n����.s�������n[I3�'B��Қ��ɥ�Ʈ7��(�iT�t��_wp�q]l��!c��L+m�T��%ٰ=��C��_=I�gQ�i11�h�U��0�F	q�����4(:�^QjǄ	�����TJ�(E�k�z�X�A0������S͢!���j��B�����<V�/rdB��gd�������ƺ�ZFdUՊҜ;�1�f���V�95 �(�t����a-p�l� ��A�e� ��@�Rh21�Yi�J1����s�:6-��E%�+
��vIT�:�C'�<>����p�$�#h?\�6�����M[�OT�L�-�1���M�>�Si/Ɏ7�O��	2�W�]�1��uhr�0B�_������S�Z_�Z�/KI�B���J������w��"�͏<���t���@���Fy��6����2
ԫ8�������*U��n�Xz�07��hB�E鏿����B���z^(������ẅ��� ��Pc�5ʣFC
��@\���">�'7+�A�F ��H��[X9fP��wi�6���
E����!��=�{ �?eB����s��Y)nG\.��S������Iy�fUk�)4���7��uq5<N���~����u���Ic�{+N�&V�~�?˄�gQ1�@G�T�WgMM�ݏ[Y��ԫ)�}ς����\�7��`'�4)g�����89���[ڊ�R<h� �7��)?�R ��?���}	�V���2���f�n%VyD|�px|��b�Y�����-�lp�����x���7�5^��j�ߥ�a�A���M�%��um}��F�qS0f����L`n���e���_,֮�eP�����c1���?�tS�O=u�+7kiu��(���J����qv�%W�Oo��1N��408���i�5Q��ӄc)�x��v�[1��=���@�$��I�ݻ�X����S@i�26����������ka��Ffrŵgx�F0�Xf�S��7n�.�?z8�t���f�� �ū�7���/0+�~�	�6!a�-	��}�v�S��ՙ��f����D'\5h�l�h�w�F���]�P�7�Zi��Rd�UpYt"��K�? ����G�Q��)gZbEmW�H8(�Лd��*J��4�[�M�Y��~^FA)��v'!�,��ʠG���#�N=��\�y�40GlZI&7�fM�b��<)9��ğ,�~���n�ǓJ��(N���-�{���3��>�X]����~B�t����Kf@tWA�����s�Ӧ�0��fE iy�9�c}�H!�/�<Ԝq��M�ur��N�u���S�i� �B�Ka�{#�im�- �Dnnn���]ލƱ�5�n��Ⲃ���Ydyf*N����~���m�����71���7�1":����S�����!y���g�Β4I�]]O��������h3.MH���7���``���p���q{%v�}���C�����x��-����K~�8n��'��{{���B�Mחƿ�'�C'T��4'�f+���#.M{�z��HL~)���&-z��};\�Pa�0f{s̡^S�]�3�i�ܚ��=S����:�Ês�V��&ܧ0(6��A���5�m�b�!�ńM5k�l1��ݷr����죙?^՘F�. p=j���L��y��@���h`�%4WpPǒ�EDE�?��=�W�}�������@Zt�c3�t�3�ʸc�8�2+?�M8^���\3�ZC�!&�� �.�/wc�Ԙ�X�my1	�h��茀�Ff^b��5�~m���J���(��J�,�6��fΈ@��<�wr��7!122�͂[��N~t�}	a��͢eȦ���:v���+�qv4�
>Pp����ӳ�!ཌྷ~6��
�&NԻ}v�c|q�$�� �Ấk!xaO0�(B�E?pc�_?gx�λ�}pb�:~z������Q"�G��Eq�ݮ�����s����	+"����yڧ��x�w�C�E
4� |d��tR8��R2��b�MB�ˣ5K�Cg�S�ǢX,<NRs�y�kHH �_����iz^Ļ���LH[�)���!�1e��<���>{��Pq���>��M�i�(�e��s8�Э	a���x�Oͬ�tH�vbi�n+`2��'ʛb��@?�Yl~�\�N��l�iM�2��8o@�.�=�o��+�F8Z��+4�>����7��I�h-(�>ǃ�Ң`E�$B�����/)���2 �Z��*^� ���Zf`���P���1���ٍH��!i�IhA�/x�`��p��N��Y���~�Ў��Wen�o��~#hOҘ�m?�5�������><0��R��6���^��ʱ4��}+;~=�ߩ���M�W���(K��ݎ���U�e�+<�:�V+iF��d6ë�A�p��[� M,������@Ԅ��`���*g*Uײxvͥ5JT��
&�2��]@�8=X��Ц��A�;$���kY�����B���,V���� |VN��/�/r�G�Xʜ�֣���ᣠ|#a`ˁ�O���9i��@�&��ԧT<���A1D>i�-�:�>ؕQV�I�fxZfQ��h>��?��bx
Hj�D>'8����َ�5��%��]�s�^|�����"��p��u����:��}�v�������وJ�t�c�@�a�k��4��K�%"�l�02* ���K�AI�^�k�M��PL��2^���	�|R`X��`���i^�g� ���19X='���76�< ��9RF� ���{��^^�F�e��o-��_��xh��_�7�`f�gkV^s{��y��+�ى>61������kn����L��Md|�}+�!�g��;�&�{��)H �p�v�&`�����A4,��x��~d�mnӂ�*\�Dܺ;Wr2I�-� ���c`7��X�%�f�RrV=��&
������BP�������ae`T�:ܠ��Ŵ������6
������m��+}��@8L��������o���ll���@aHqёK�P O��|e><�L�����?�����8i�h�w���.��e�����0�� "�N5Z�ɏ 5�Iձ���$�C���մ�:n'���RU���
�ӟ�v`��y�������}BQ�m%>D�� ���8���_��rà<�*SO��b ˂M/��h�1�q{��>��<\�je���N��^I���wssl�:�3���IoߏG�%�N2�.9`db����vmO�\G
w��dZ��٫P��ЙU�6p"]|���~<��ld�
w(�'����K����E�Ȳ�v۳b�&���I^HJR����JJJX��55��H��Nk��m����2]>E2?�]BB¨���B�c,|����M�\�nnf��ot���$/YX4��$��\22����c�L|w�S�ϐ��o�����#�� �F^O"HFR��	bmN���'�����6�n|yPq���`1���BEur^K�(S[u��͛bI�|�;I�m5��%up��Ʈ�A�)S��'��X:t��׊������Rᕑ64�T�8��������{�F��n �[��G1Н�O�Z�|�ɯ%ʄoj�h�
�q��8�
���������UDn����]/��1mdDW>����˯	��%΍J�e]GKu!D$�v� ����n�΍(�ɕ���wxu�T��f��Jhk��^k��!�?$��H�����T^�.�S�J<���Y�����E��-G�!�ъ�{C�mhL�=
�d�1mj�)��~��~˿)
���R_TM���Fu���m���ڠ��UYv��kJ'>�_F���v��zW��ȟ�EFE5�z�9-��}+r�z��Y�/�n�V���Q�U��~�� ���t���LW ,��3V�.C�!l��K�9l�Ym���C;�;�Rm�k������7��>Q��6'NY�}��Y�Q�]���p�z�_RZ��r¿$��鵞cy;i��ӆm}"����u��3�6��ҋ����	���𤗕'��@J:T%U��:�JR�{�!Dċ`����W�w�뫙���c�=�K)�F1%OQ$� �*3�K��%���
��o���u��F�߷�t�w��5Q��6��n�����FlDAa��9�YMg�縥
H��ں:��G~?�W�:W�1]ߪxCj߾U�0�!Y�ui��Kk�Y~�d��׋�O���Mҫ�G���/��������`��-���ǐ��[XS�u�� @I�:����5�[���1�iU�5^��''U�Ǟ�\��ԎN�[��7+ೋ�-�߸%U'g��M���Ã�����fm��@���d���)vqo���m���`?w{/��Eժ��O��@
�m!���,��!┡��4�̗�������g�ȿk�.-)�$*;}��_m;RQ��|=� ��������ǎ$���v�^����؀ ,}��n#E�2\�t ��gQr	!u���Cg�|d7�*� q��jL$������-�ӓ�}:Gʌ�������&��(�}*ʰw�M��?x��J��f�/�ځ:~?��e�=T�{��6��:��+&v'��/���͇�M�o� ;�|��1�ݿ!T1�P�k��V9 ���'%���G��}�#��t���b��%�k*�s��rsY�fB�:$%��f?L��̚��#���4F��/\#�V��gG���ݙe33U��Y3�fst�E���W�o�kF%K�kFW�f���^@ڌ�N�����ˑ�b�7Cl ����
X��å�[U��h�~���hS�>�k�ۈ^��)��)�7ܟ5|!4��fS�����}�i��*5VTӨ��@�ٝ�"��˼q����q���BV8�w�L|sv1!N�籸�4��\�/��?��<���ƾ$ʖu�-![�Q)J��!Cd7#*[RJ�ɒ%{��/�KY��kvf��1~��y��y�����s�9˽\����}�?;̝�|u����'��'���'��k�ҳ,>
�l^EW��Ϳ�,������Q���t�2۟��) ��Rd��\i�,���/f��*�$<<���GN�Z���VO�I��ח���W���V��%)�.-����Wz��"���2G�䃨9�'�`���y�}B'+&�ƃ�?��.��hk��7�}��KZ��L�j��H���b>P���h���y����u)?"��i�	��vz���
������/t�Imɘ�l��Е<b�t���S��ޖ5����Ę���_KCp������ѯ;��ӓ�<�Д�q_^���>c��lӑ��ȢV���V�k)�U�̶�p)�t5COMU�^ʂ�:>b�Z������6�wj.�̬�p�w��مU c�_	��C��X����犿'2�tȢ�"�O�����$O�90a��]�]1�u��P���\�
�*���i��K��I($���ˤְ��zB����D������b��R[	�us�ߒ��~�NvJDIPuʴ�饞��oN�U0��>�Ut��)o��%�j�f���_ڥ�a�h+�!qw}6���,ǲ�x�s1���JLdu ��:}�����X�z �c ���b�ͮ����ܚ��H�y�]�'�S��7����[1p���GGG���ϝ�� B���s�����%y��4��`I*$|÷}p#���x� ת�˿iy:���	��-���� 	�����;�13�����T�=�K�����=,�U�d�ۅA	����8���s������?\�Nyd�@-�x�����R���ċ�J�Z("/Q�j>���h ���0¢A]�v� �� W����\g��)��=���ݟ^5�I���:�uyd=�]v0���D�8qw#�,.:}
ມ�t�w��>��t iR(1�Ë+�!� u�Ώ{�xd�&��������a��4�9'&�.{iɕL�E�h������ҳ��W�$[�S�-�����
K����}�;��FN�쏮�����F��k��=M��	' lV�^�2�3:1Qu�븙��T��x��T�zxkn^A���-2|�~G�Q��o�$���"���/_��;w�%�z�C��|XKSڗ�-�L�
�w�Iv���������>�H �����]s��ǔ�g������傿ezr���MK�X��O`i|ym�OU���\xJJJ�At�KI�_�qtr���"kv�k:���ɪ���3њ/�\�(>��:��aEC}�z�'-�yW����II1c���6�2D��hO��[j*�8����n��0��(~|��`xp���<���P��8�H�g�ɟp��)���&+܊F֪
�"q�������Uc��q��#��p�ZT���0��/s���;jLv��y�N�X���m���o=��i�����&������!����=R�l[4~��"W��"8�^�(��>�l��íyU}{�P*�y�3����L��Ê��_-±�1��@�o��Oy�:J&tv�`%�v�#��ɳ��(�ەi��H>�n�P���/�15c�v_�ȑOѵΓ`����u��B�^1:nld����lIjJA^�[zέ8��RJ'��cG�<ñz��[��c���/��W�q�kV'G�����
�y�����{��ܝ;���YS:�_6y�`�ړ�[����&�=�1M��Q�W�x�͖�O���O��^0A�����	r@l ��68�#����bk� O���Q���;�fCΪ��GW0%���{�?�z���QJ%���u���;"��_��}�O��٨8*���G����0�Jҳ��C���ѩ�W�������5�QvI7���a�B��9X\�U8����ޤ�����l��;��b�ep%X`�\l_eQ�ZY�Ћ��w��cs�P��?��7z����V��Z;��)v>���~��6���6��Omb�]�#�Y�����b��=��[a^�U޳n��q�E�u$Lbe�	925ݤW ����~u^�:�x�G� k��<*��IiD���8*'g���J��lt�[�輯���ˇߴc�0o_7_�VT<�W6ŰҤ
*7qm`*-�"�H��zŢ����.��C�~/���?��l �8A9�z�9zl�N|���}g�y��;Z����~����T��)�5����k5;I�S-�J�-Ku�|>	7�\~F\g[��L��4ӎ!T�q��ǵX ��&��F"1o��}���[E���c�?���M��TPs���tQo��I�>�W��#;ߨ��+���re+����b�ѳ��P_y�oـ"o�ҋX�S~���@�����^�0�x2�%�����&+h��U[��֐�o��2�E�Mq������ϟ�����NȺ�g�7
9�7a|��z���J:���Ј���a�-0�`eD���$*�yע�9�ߢ98\di[-9}��A-�o�M��[0q�j2(S3
4�����k��gP93�F�>K:��In��Ƥ��L�>(]兣TV�Q�lpI~��
/5K��B�ptB�3Vr�����m��/�8Q3C>bծe���Oܺ���De��j=��о�Ru��s;��v�+���ۭ�:�+8�}��0���D2+��QZ<�@��M���]�ˍ;J���*���Ė0�4�)��,NgA��M����4����y�۷�����9\����3AR���u�D�\ 8�*+b��(;�{�4p6�(V	��h��]m��j�-m��7��u�+Z��%�ˢ����ۧQ�'�+°,P��]�pOz�����4�9O�l��/) #?��1���d�dl��>��TW�~�HP�y<�a'<s뎕�8�9�3sSSS�x�Վ�\����QC
l�ڃ/�M ��	���p�L��{���u�0H�{�����4�y�N/l�ND��Wɷ�K���:,ך`l7ܦ�ޒî.֤WE��I`͇t�+)�>ü��@������e���e�^�x�Q8֛:*oJd�l1p�p�k���TFU�]	��[JE�߱{BgE�Σede��ɞV�L'�`ʳp
�^!ň�����3�RU( /R����}��(ۡ"���w�.ܟ��lǴ����������=C�ϟ?7��.�N�&��O��,Fi=� ����*��������S�uF��	(�瘓���O  ���m�6ǚb��#�����;�6v��M j�(�Q����@��e�.�C��iv��jb���p��'����ߥjٴϛ}����(��3tW��m����.I\���ݯm��ע�{F���U����̊�lG�@�vY�v�!Us���=$͡���NK�}��A7�&Mq�9{�ll�`ի��sƷ�WP��&���W���Y�w���x�����u <I��d�+�.�y�����+H����۳+%K��V~:����'�����p.yv��|�c굷��K�3���s�BW��W�yVU5a�b��+u�U�#ug��~ό1.0f�a��ʷ�G� ��J��������
aZٿ�}��
.�ui���0�
ܢ�;��3η�$O�ȧs �&;�m�Pq�2�~lt���T�Xԡ�]%�u�������+W��cc���wvE�&�یL����XJPvp^oyǷ�'��I�@_�2���Npɀt�4�=8�]�� 	J����W�`�n�Q��ο�����Xb�C��w�6e�v��3)�|:R�t[�f�Z���T�y��\�* ���j�ڷ�?�䷪4p�S�`^�t����m<�a��/��03//Ҝ���	�
��wl_�m}�����\�u!pf)n>d�n;���B��X-����	 ���5prJ��ԣ�4����CVx�CJC>���H��I�6n \���9]����	��(����v�̛��jH�G1��E,����U7溟��'��$p��۹��dѷ�ch8��.�_�]�lh[�<B��m{*Fm�p���)+3Sk�(�NN��h������ώj�`u4��K�7�W��C;7�%����0+��J�#����|,4.����h�P�po+�	�n��3"C��Oz5m�y�T�|����G���b7G�v�^��q=���Hy��~�W�ȣ	:^fq�<���A��3����">�_[[���C�y�M�c����E�m��6��B�q�պ�<�#<o������ۘ��]�_�n��	�"�|�����sk�A«���'��\�Pҍ8�+�{��з�dK�K��U� �Ȇ���FxZ��l��O��ﵡ��^�HX2MX8����7�L ]%�g HD���O�3�i��3�zd���F �
^�"����!EGk�c�j�g4�&&>��ྲ��r�g¹ׯ_��(��Up�?��Y�J��痷�y��d]H��II�0�}f��v*���uñ-VV���ɉ$�}>vP��j�[�Wϖ2�3��̃�����W�Ǽ�>�j���b2t�������d����^%��4�*wB�-ze�dj�7D��a���27r�^�.|t��k��`"�1�̜%N���W��)SL��Ρ��d��'�a���E��mx���򞤞ED��ҊN��9XAF���/n�p�:wD��\�N�n��r]�~�pؒ)�E}�C�R��e~��3��s(ע��V�V�`�� 	-v�+��0*��:fb� �h^�U�?��Y���:��������(.��9�n�H�n��J���);��@�ܻ�?����W?���K��)��;5�k-�ۗ�����qo0���%#�)��r���z��G�U�?�rX�5����<�8|:�޸�?~X㽘�qE��~mOȘ��o�n�7q2���i�������l�/4gw�!����[F?X�h�|��j�+Q�X��b�MTX�=h�����"^�٬J�
K�����RY�<�*��.�E�6�c�9���TĞ0��Oy�Bz|c���σop��Bt������ώØ�,���9���2��)3 �����u�
r,|xR����G���h�Ȣ;,b@D�om��^���eW��C�i���k��WCg0"��3^�.��ٰw۷�C��C��%�ɍ�l�"��T߯�����z�'S�x�L 5�SaZ�j��>�v��D`/����++-���|��=��x��e��ۂ3zF�~2��"zI��4�'�o�^H�!��P5�}:��̪ۙ}�cWMHT�yo��h_�h-�Tṫ�p)ы"�={D�qÙ�΁�s�	��N�f�.�%�z��*=n���o-.| FGw\��Xr�	8�6|)���P58�'ӗ��r�4���c}��$*��S&�{ok�;j7S�([ñɯu�j���P�� � ��5?۸]Ν����P�%�[���S��
��ث!�ÐK�Sf��w#��2�X0��=f����X;�?$�՚����|Ĩ�	���#�V�#�/����Y'�nM���yR� �5蛓ω�{�� ����ҁ�X�V��[��\�}�4q�d�u�h_��`]
�4�*�``
(s����/�}�?a�|�n����rW i���4�`�~xt�5��B�ԍQ�6m�������+�5�B\��]:����[p�2�X�|%CB��%��O�S8���`t��H)�+U��4��o���o�N� wW�i3;�S�O���L|s����wɬ��J�gJT�]7!�s�3'��	��GUr��y=�K�y�M�1�9���R��-=��4_E=[V�`4�AaF'�n�U��K���4����z����	}�BS��ޠ�>Z,�<[b}kM;�~}n{�������ϸ��������΍��Y�9Q�yE+N�	<���I�'6=W����Nʄ�CU%��LhrC�6j9fj��m.�JY"<�a3�IEK����`��4��r�P4�b�A���]�L�p'�0o//;p���n:�/1rHD��uFcb[���&�� $(�UMj�eBOV��L���B�S�_y�S�!��p1�(8>����	���S�������;-�_b@���Oj
�%�����Sk(��y���Z5R-�5�z��ǉ�ffAǷUx�@0swX�����#�Jt��
�����9AH�j"wb��$'C�em�?��y�B��xV��*J��q����#5WZ� ��(�t>M��Х�I!b�qu�W�����I����a`C�Q��M�f����y)��@ϩ�R<�qA�Αh����@�)ɍ�h;�SN��$QQQ��m�:�8Q		D�+��3!�1�=����5�Մ����9����Sw# "�����˄�2��r�H���=9?sCK;�*M*���"�]�Ռ���L��DQ���&U�օV&4 nA�;�o8I����0�ާTK���z+�cd ���v�$f

\3�����DNI�����S�"��-r�T��3*
vUw���U�k�e%�h����5n�Iw=�_V������L�V�	̼Cɇ���E���[8����|�svv|����w���}�M��OKܯY4&�9�d�>He�ɫ�z�!D�3C�4PC*Kj���M�����Y��B�@��2�zդf�@�v�A`�z��� i��5�4�!�=2ݎ�[��!��.�JW��[J���zX5�8���6	�=�>s�_^Ƅ,�	���)I�V}��`>�-�>V	բ"�R	���rB`-R+���V��h���h.����1Z����h潁Nk?\);�>N�e�������hhh�k�Iiw��a��Z��2�QeW������:L?��GH.Q5+dD=�н@x¨��������{K��B-�t�m�%'�U�,v���Nq��LjnJNt���l�XZ�c�K������#�q�la���CĐ�"��]%�)�"��8��?2g����2������U.�����[�ۈ���}*7,4n��>X��Q��T&J�<�≷M'z����!�X�kV����7�����H��:�(���l�Ok�a�����A��Z��m/(Q�S�;����;���;&r׵A7�%�/��:{�-~q��}\�a�P���0Ne�GV�h��+�O�|��\[U99��V��y�#}0/ަ�ˍ2u¹�#!M3Β
��y��\*��Jk6��y�����?	��	u<�oEԢN�Η��_j��O#�b������)�Dp>W����?����v�����
(z�)���1����� �����.ww��h"�YVzv�4��גKZ<�0�M�ԏMm����ۜ:��f l\X���DU��1Ohh\����>���4�w��>�!�7��������r�5�.������@�;<x 7����M/r�9�<�!�<�HS[r����)/��{�)�66��/-����*��a��L ��yM��%����a
�a�x[V��DA"���YVr��he�:�ŝw�'�=a��ݎ��W�OZ��!}���?�o�ܟ���H��Hi���/{���s���B��y����c�F����K�9�U��QAA�U�l@5RaP���� �j� �w�r�n��@��P�C�\��^��f��C��.�*�S�Z �=	*"�f1��Ǐ`X���h�~�\�?�%ka��C����I�I[�>�|�z{����3f�
�ߍ/ǡ��@�p.�)��V��d�b>s�=sQ����~�*wrUT�`QH��2ͯt��x���}���-u[K������J����ޫ�0W2/O_��?��)e5s���%�,�]=�=�L͛���~�2σK��_ޭ߿ך��ՙ��� �k�Q�`1O�V��^����?(�۳��_䂣��0�O3�`�8'�T���@(�6frr�	���"A�`�=��g<	p���\:9Pc�B[Z�}�({#cEԀ�N�bҡ7�P��,��/i�����7���L�oN�����5
mAXٹ�9��C���J��ր��M���]G,={���͇��W#fp����P[���_]1��Zfvvj�wt�ԲM�����e}��Ɵe�}�����}��VȌ\���bk�O=xL�	�mV��6�+(�H$��[�u�=����A=K܇�a����.�$7�e^�����_���4�{�,p.��}�i^��S�x}M���}�����J��6�U���{�{-�s�cY�����o�T�4����k�wD����:�N����1�LTn�V��7� �&cB�����7�:,\ ���=ѣ��o�CrC�`�S'�0��͜h�2��]��Ӓ�����]$��z(%��¯rk��,�%����('���Ǫ|$×��B��펄�e�5���'&c�͢*����a�'0������2���@a���0�?��6�$���I��AФj�f���=��Ɲ4Y���� ��:�P���D��AH������k/i����-~�{����ճ(uNf�<�+l>X-�-j�"2c�k�m:�q^?���di��S���g&j�l�څ��PjLb�.����K���]�Xk��<���0���D������U�K�+�?�5�	Pf���NŨ9�_fV�da�Wy�V��\ �T���Q��в�|���c�-��/0���0�۷U�XyO.��k�F!����r���*wV�V[ه�D��m-͙�:W��+ѩ���8��'�ç�G��DA�Q���f``����>������4�=��ƌ���<�3^��q��Z��:L�UD�u-eW?Մ���w��FK=�g�>�J��Ӻ���%S��v�/��U�����\�jG�;�%���c�\�ٸ�=�iZ��灠��	�v�����'��a��N��!�Xcx�Mm�Kgo�k�'&0�'@,1]��R5����e��|dg���C���N'T�WX�%�g,2��gk������sg�#K��-��Z�V���B����=RF��>9h�8�*{'���Z@���mD��n>"�@�D�r�5�偐h������i.��������~�̔�C��'�8:����QK�n)x�_K������Hœ��O��k
{z������?i��\o���4�ٱe��Q__�/��X�!�(s������2��zFTH��1z�z�vU�e�}e��S��'*����&֨ݳ��'C�ڡ��psCSgydHj������Ѡܝ�w��OU�k�t�Ί0p�{F�ܘ�Ep1����m��^)�`\���'��lM���0�}4�+·���+w*����*;s��Y&ם�ǗX��Ĕ����D�<��+Q.��B͓�����wb�թ�
$�v �B�y^��3+v������6[�}g�>5uo퐌�Ɨ��E��#�����/��o)�v���/���"+�V��WN�3��.�	}�|�X�/k�s�'Z~����Z!,�d�C꧈� ���ܲ������٢t������AJ�˗�:I*��D���b����̴�ƌڸׯ���$~�Bq\���B�qqF���C!���*�Ŭ����3��^B2��@6<���@�$s~�����[�����[�Y)�j��7������<VG�V��SflC'0jP��\� �0�-���yW)��B�BI�p:�d@���(�OL;�qޏn��] /�^me�$5-M�s^��Ųi��u�S����̳�aH��Q��͂����vvv��ȸ}�)��$��������X)k]��	�V^Tr���ܻ�ec�nAֿZP1���f�_�X:?�lv-C;�<��?�Q@+�h�%v^Xx�÷Yϱ�QSuZ�X����h3}�߁�QHۧ ���׬g��T�y���~��^�~���1��EeZDFtl�\�(�Bx�@"K�a$���d����Q#��1��!��Ã�ܱ�����$?��{m�lcd���O��P��9�%�/�سb��{�	'(Wi�/�>ػh{�B�hå���35�)�É��!:�F��{zz���k~�uW��J �E_��K��d|��C��Y���f�d�� �D�f�lh<��s&A}���e�g�/`�)т/;�/50�0opJ\�7��M�a��<�6Ã�v���b�I*�q<��g٤#Iu!�k��eJs��9A�;�``�to{��K*8So���D�O������&YZ�5p.���+b��Sz|��T�S�����Z���*ޅ�[���r������no�gu�0C���o��y5ҩk۬��d"^��Oz���Wc��ZTb��x[m�7Q~�e�2��4O���p��f���.�����v�,cR���S�Z�vLe��2�}�A�Q�I��Kb�����+83�� **���q�Y�Y��L8�Ï�g;/̾�W�cd���]V*�)���"�jJp_\��#��|�hU�+���B}/��k��rw�jg"ۼA���T��Qۖ�}�	���4'�� ��b�Q�=
��Y����x�� ������]�Ir��O�#eџ��_a���_v~��Ѫ��������g�Bz�DK�(mX�y"����Y��ƥC�ޅ���q��`����ޛ>���Q�kѠ�I��sl�nO�4��R���Ë�����\:w���f�$�@߭�Or��{��)�L�l�lB��^1�@�:̪8*�+w�霫3��+�kf�G�b�������F�-�P6"��~?��˗/��iq⢎�
�����
`��H~1*���s�c~k���_B8�_��5�P�t�
n?%�>��y|�ǒw��)5�����U�YGNR&����E���ơy�]{�ȱ/���}�rq�!�v�*����@��Y9@M�ׄY���� �i;���o���'6�aQ{E������.o��Og>���y�׿4����(���ڗ�
�,��1�X�k�2�p�W�TM'�,��=߱Vf���Y���&gkF:2���8�����ozF�.��� �ϫ`��ӹ�5Ҳ���t}Tԇ�%�tO��o1,"�Q���˖��3���!D���)w�<걓!~u��,E�M��&��̓�������������j�***z8R�ֽs��,S�&�Zk^t3�oA|צ���Ԛ�5�m�Q�X:u�:L�3�@��	O%�TvnLu�#��� ���mu!N2���c☶��w��a$����	�J<v[%��8��x���]����3�s�#(�5�hJ�����I�C*J]j'R��)�<�wt�bT_I5L�X��{�ߋ��+�����[Iٶ:Zi�߰�$Y�J��ɽ��Q&2?٣�ni{���Y�Ł�D��ۦ�!�v��̐��pcH�
�%Oz�Fw�:J�8I�.���4������Qa̱��QC�Sz��mc���Y�?��ٷ��C�X���j¥Q�'��İ>�-Τ��&��/�<gD�!�S6t`n�{�f$�B�k0�j�v}�S�\,�%�ֹ���0%����(]t��}�^`�����aѓMM��萫_�<6m�=�R�p��/�'+)����v�QbxV:�h���xڹţ��UO �FA��B1��>����9��ӗ�IT�bz�?����K�hH�9���0ٸ���g0 x�` N����;�K�'�6�BS��}A�������&rʙ*�������0�����5��*m�A�����i�)��/���*����U���!
�%ۑ]�E�w�?7${Pw���Մ��� {K�0�|�-�wݷ!�Y�}nw����D�{x�RHp��7X@l{Qwj�+��pq�K���-���ѧy��c���Py���۾�׀~X�W�1� �t�o�e`��������HhK�a`A��~+G�&+�s{��5�l:ȅ��(��",ly�u�����k�Aq,Ӆ��9H�'ԝ�xwS_�K�&�����ˇ?����lcx+\aA��«��A*�N����v�XVy���	�@"?��*����M�t�:��1�BCu�o.@��l�S�L\g�5ts!{��zͮ�.��Naf�l)T�58��	�q�0w�x�Y�NŹQ|FY���<8�Y���Y�����;��������(���u^Cu?-ɢ��@Xx������h�'��h��j]#�=�ìAG��ru��1�M�w��i֐� P�|�&V��� �e�V/8�Q���Q2�Q����� � �c]�i�[bw�<�$�"�i>D�uf0W]I��喭pY�c�s-�d�o����A��vr�պ
�����:�d��I���!�x���ݲD�z5����ŁȌE&���g�sP8�:���������"A#�e3&g��� �7�%;�$sw��	;R��[���]Y���X����W��JϺo��I�������
������E.��!���Q����i##w?[�|�y�9	�O��*J���#^3�/��R����� �|m�k)N��UO���N�b�S_����(T��D������b�,^�Ws����i��&� o�1=7����_AԌ��Cܧ�N	�z��n��G��e-M��4�)~�Io��/�ggg9�N�3L�6C�sr$l�뚘	�"E����Y�[b7E[�>!K.l<^(�S��o�X�W|�`o������c9�|9�C>����Dm\tb�}���� "o����M�M�jM0�'h�@$���}3FD/��G���Vh�r�f��)��R������<���!�Џ߱]/$���N�r��u��i�'.�}��8م�Z�ǔӛ�oŋ����u�\��pttt�c�s\a��C��Ի�]ɩS-*�c_���'�� ��7��"p���P��d���F�P���@�� ��^���3y�-�������lUB�`��O�,�]��$6�o�{�,F&��f\_����� ���v5�������+�,95
�<��:s�&r�ٳ�ᤀ��)�~,���d���)y�)���[v
l2=����i��������nx� � ��1?�ف��G)K��NR�Ic�"'��و�8��������@����0\�&ɞ�S�a9�'4*�@Z��G�ZS�!s�XJ���W̾��KO��I�<���
��~���֩�
=���ߍ\���4�qׂK`�K
��𼢥I���w�c�\�W&���n��̗�V0��T��5��3|�8��x 2D $?1��R��yK7��U�;A��n����S�/^�K�'�t�J'iW
�z�9?�e�]��h����燅jr?\.�4�LY��;K⳺KB޺q�؆��CsZ00d�ќ����/+�����G���c���7�پ~Z݅�I<�L�@�ƣ|�D#��2]5��x���.�)�zk�-�z�68][��7~�4���I�( ��!�4|j�F� �1l^}R��� C ��5��ߐ8�^jD�jii�U�uO�^f���r�u�� v-�q�9��cD����J/�%�)����M�=����X�f'�JcH������6��ZXٔ;�Z�	�?�Å�d��p�杤���o���B��M�-rn�ފ`$�R'����Q�8̿f�귝�����;��~�e}�{�чe���@�[����3~hӟI����
w��-��rU�;��T}߀�|�.R 5�0k��q���̥gu)���ך8�=F��kIה _�	�/r�+|6һ��j��i�]�D�L�<��6NU�M��Czz4�<<.Vo�Y��}�����Λ�'&?����
�h���.�>+��#��X���v�������ѭ��Q��Ar�߄hc#.�^�&��:Q���빹Il�PhF���TJ+[M��Bۖ�G�/v��o�~�3�kH�soh S�𬬬 2ڮ.&����8����/�qr:�|D:ɘ�.���B�#�	A_Ȣ$P���V�|�2$lB����߿�f_9���t4�������Ս�� �R��PFTWUS�`�bQ���R[�|*%�+j�AJ�i��R?9�V�	��T;0c'Z���h�k����O�=e;�� ax�0�|��Zס��L�����>�%@����b�R���!�y�pN�Ć�s�^��&UZ�W���:�G�G	ø�`Z�W�6�4G�S���} l����l��������e~Ḡ���
�����
ѱ�E�)&��"/����� T8���:C4��'C8��cT(�w��ѵ4��`vR�qug?ec|���΄�YCݎ�1��@���9-|��o��� �s'4���s�f�VH(_>��M���ؤ��C} BS�]j�J.(88\A��3�ɴrgMt��[}�<�7���>�����ş���o.L�M����ZY l,+���y����+���P�����w�4���r��hp"�"Z!]�}F�$��/2�T_ �Jqċ��W��՚���rzsZ�hÏz�GY���� �N��|��T�&����`���<j*k�.[t_ap?�܅�ՠM"2i3˾l�'�.�Rl!滬�O�jv�*���i���KJJJ������C|����k��#"I�1 �3_1�@֓D��zB�Ł��V��ꓚr��I�dA݁��'0��G,�y:�U|��'lT8�'Ʝ��� ��/s����a0$={�bO����i��Snaz��<h�x54r��K��>g421є�o���T0�WtOW#j�33[�~� �K��{��*?/�����3�M2�Τ�'`���k�1�5a�,@���]���$�c� �1�5��QJ��4�o���`�	!��Q�J���U-��By�� �퍒Gh)^�R�����{�'!��(�$�Љ@�zL"x�~�L��$~\=g�y�J=�wI���n%�X
0"�P̣�4ّ|5䜊������5�2^�2<xw��`�|�Z�����(�x��Қ�~{�B>v��b��}D������֚gE�j7o@E��z��r@�*c��E�|�*·L1�e���M ��;���A�@�x��)���1�IlpЙ�P��'z�9I6�(B���W��Mm�O���<
?{� 'sѷ:=���Up�|��^����R���j�3����5�Q;wt/q�f�@��}WO�z��B�e*���J�!xAF u �s�\�΀H:�z�W�2dKW�07�bZ��M���&����i�ϥ���8�a����Z,�`���[�m'-55N��ϟ����kU1V>��+���|��w%��K�['��1��d��7��<xнC�)��/^�l����`3��ݿ�j+��Q�&5�@/��u�%�0**Oh�HNh4��/&��8��EҀ�Q�Ph��.����P�@~Ũx��	/hK�G�y�F�D�~&*�1�]�C�V�̌]>��t��}���'�M_җ^$�k?b �+��G��;�A�a��F����տ���ex�h���p)�r�G{���(=��ʯ�@�S���߁�2�������2���dt��P�ݒG@�m�9�˾2�Tm�$c�^Ȉ2�[�k~D��-���EN���� �gk9��sWa��p�Xo�	n_J^=&��|!�}��NZ��w��x�I���@H������?:���w{��vP��٢xͧ��y3JK�\���e�YۭK�kN �[]��q�~�n
;
24WDt
F���l�I�UT���X��_��`�1����^DLfx.q�L����ά�.���w%&`�ϒ
z!��?;9P�.L��&g�f%6��x���;7��EHwku��ʰ���3�rc#9�}�y�7HC�@�\�<��+�����37�>��P��h{�	�ZJb�ˑQ<ƭ��=�}�a'��7`�& �<ԅ��{���ׯC<���#�y;�_�Ek�'O�`�Ǚ�����v�F�˓$9竒�g/�o1lQ���bu�K�$�,�����g��
����u5��m?����}PTB$���e����4���Ō�r%<�@�?U���ll���"�S�׮�@��֢k�
R5���S���_y��ܪ������1 8Z�<����b�O��r���4�m0�����L	��/���pSB*?�T�'W�=��m��L�)�<��/ ���l#u�~i�x��F3�N&�@�[�E�Y���'����	����m0a�X���zlZ�3��/;�i��{���G.��T�?Ow?���"��K�3�-Nť���	P�|cܳqś��Cۏ�����{G���p����l� �{���B���/\G)�0E��Q�����ua5�/,*)!qA�ĥhW�+}N���Җ�}���W�.OdP��W>�u�r���;�eQ$3B��9YT�ej���Dz���Ң1Rj�{�.��7Ѝ�h��E�3Q����*�E����:,`@A�RwT�Tϱ�����
�����Ձ@��h��������dL0O��޼y#e����I~����d6^�,#��� ���
���X��[�gK��;^�(d�|���,�@?�vb��N�������U�6}=q��������kǫx�,�������ߪ�J1!��t[1�Cc^?�u���Ԕݼ*�P��/�K���l^J�1�lcGj��Ph��s�%!�I��f#���&$j�'_��0�� ��aLq ڵ.�>>>lllv*-s�hbp���.�����:��]��"�N��=��>Hf��d�L�yy
и��W*��I�	���W-�m|Jw-�qJ�x�,�t��=O4`k�;&�� I|�{�F2�1M�#�(d�������r��'���jQ	��L4��>�p����1|C@�,�޽{g񛼿�P�3�R�b{}��cZ�Z>ǏQ��"�tmθl�pH�m���i=� �̌�s�x!պ���,=(��������������vk�����H8��o{��ګ@x�n�����/ϿRh����/�r�F���p�$_�k{;@4��B�o#��ң�^���M�_��B/��d��(�u���Ƀφ���`e�:�wW�A�l�t�E�Z �c%1�o[�?�_�?~�w�C��!�Z=�54V�W�*ce��p�Y��w�벲@�cw�x�F����DJk�}S<O.��d^�^��6�Y<&� �@#1
�q��u���l"|�__���T���y �{�?���$1JH�QD����I*I)	W�dK�mF-�B�)KD�fߕ�e,ٷ����`�������|~�fy���<�}��߯s�c��E5��s�����4�:�k����^a4����zT`o��F�Қ?g"
Z�s�������Uh�Մj�s\�?P��	"���S0Ƕ�D���m�y1`���>�F��~l�l@4t���ׯ�r�ee��}HM���C;~��iof���y�}�{���jCt��d��f������p�f�o:�ε���:)�ѯI�����)��F��˗������byn8��7�?�x�<]]�e���vF�w�� Ȯ2�%k�ѸC�L(\���i���_U=�[ꍢ��i�3���E.?{>�L�͕��WUW'�G��kN�QO� �J�M�=�c��?�Q�
b��.�)D�*e��}0im�뭲�^�ݻ��
�mVf�]t�	{�C�T6=�#��b�m�@��8�y}#.\J�(������tZ��8�}ԡ�c��z���ֻ�]Yg���9^�+�ԕG�������1�e�Q�+uQu�n�[���ԃh)L��TQ����BC�IRG�dkS���}8�)���/��|���VK�F�}�M���?~�I�y���j���<���%�Ç-SvI�U/y�0⊊T;�tpo07�H_ڷ����}>��u����;��JDg�zp���\>>8��	�1�2����C�2F��y��.}Ա�����`�*��U��V�IG(���7�،H$��y���5핽�{v-��V8��#��y�?O��C�ﳂ���fqd�?O�O~�J�Vݜ٧�j\�C��C���(C�D�ÁW11�gz��7����r7�̏��	k̻}�vs�%a�1J����r�I~Ӽ���G�p��//d㐿�a�]-(ɥ��8W�ʂ�]<ꀝ��Ht���9���@�2�W��Ӗ��R�y�������7Ou�5�\:M�3�z�&���δ8���[r���m�G�:�+�|s�S��B�1�̤����X&R�a�l���c]K���߿_��\~m�x�p[C������Mt�/R��ƹ���{�Jᗍ���	�'��rᲹ�]`lB����Ab]�t��[��f<���\i�X���T�b������x�|��Z���K�v� RyF\�3�_;� U[��WO�i�n���s~��]�l[f��}���Z�3�O3�5�"W��LL��@���猡U�ʤn�pĉ�v,��J~���hV�,�n�%�wu	 }�c ���u˘DV�_�}NI!�������E_���šw~�����ae)�K�$b���ͮ����.��CQ�٬#O6�W�w�85v
�.抷��V�}�7� ]�Rϵ$p�fr���گ,�������E�<��_�m�<r�-'IIH�RX��0��Qn���92�� I?|��fs�,�7ױ�������y�Č����(��y��^XʩV������hd��C����N���˘���;\��̴��KJJjal��O��p;''DZzQ�-s.h�_l��A�u����oHAe�� ��F�B�E�+p���1v��*$'hjùA�����$'&~eCE+�g�Z<)�Z4M�d�}oG���k�/�F�����k�9��/�pXg.���{���|��{�Ƀ�A�x�Y�)Ni*�h6�@�q|�ũs�5���.�'q��	�Xq���mIz�����f�Nߕ~k;^QQ9�r���V)D��G��� ���3	�K ��cU�-�Gxz�}du)g�H�t?"�U�70x���gKm��m3���=���ɕu��/!2X���($��)84����)�����e`U������4�Ik���ho&F���d
D��0gA�R�fx�A|ڈ����Q*����B�EWUU�577�X|��xt�=-�No�>�s���5k���P�:aBԗWϛ����ͨ�q�w|���nD�8v,9��]N�,{��-F{s�5-��x�YHȗ>�r��ƚ�]�zY�����*���E��s�_�� e�L��|����{����=UVRR
1���m��vv.��r9�U��*E��Fq�
%_��qbĨ����V��ҠF)n��D�����ׁ�t�Cᡠ���үgŷ$v�ڴ\t�y��qat۔{x���<r����3�T�' ���M3�Z�غQNE�$n��/pPN1�v=(X�����ɹ�<��줓�pK�8&x��/. ��垹�K��)�d��h}����t���	+��ay^e��x��y;�$Ҏo���uh�{���.�y�����,7\�L.i�"��}d|5��dg~� ]�;ꃑ�sĮ,�	Ц�\��m�v�'�,L�!B>92rN�ڕ+�E}�eCb5��ʒn�Wi�7�EG�M�'~A��+���'prtjuu���V����{�����iD�k;�r�,e�  � ��6T���!.��#s����@��fo⽫_8�U�q>4���a��k�/r�=��zv�e(�M����y�'7Z�͉X`c�^�/��j��&6K���g��� 6��M*9οE�n{�U9��Ӹ;TVa��*6@�����V�Nc	��*B�`v�8R�tM^R&D�xqb�����m"��䩺h�+Spʫkm��;2y��m��L�Z��?�e�Y�����Y�c��l�N�42�p�^ �)m�����	��'?�V�S,��kR=Fmh#�T^���c�i
���(�R5�-M��C���=$�5fu^xb�0��<�+���V���"dC ��z�P���P�0V��M!���Rv&K��ϗ�h0���#���^�:�j�	�C����gS��3~(E�8�P��RgO.*]~�YZ�t��N�G/ҷ&WrӜB���a��`��zn_p���R�D�#���8:�<�)��\<�6���R�;�:vM���x>R3D�����~wik?���s�g�����~n�]CY�`p�0�Y�Q�^���K= e1 6�P�FX(d$n�W,�vޏ���bw���5��f���=KT?N[�9C"4�+�#Ԇ��c5B��fLcp��ㆀ�;P���R�t\U�X!v�b���j�(k��5^6D��D���<����gz+h6��~ h�Z�Ї�Wf�.�k�X�;����{���M��&������g�JB})J�ugs�;��a;@�N:�.x4n��iCZGHA@���#�g�7��9Ϲ��vRx	C[J3be�J�D���0�q��
\��C)y�B��rӀ������}g�hd�� TNrNB3k�z>�o\o3w[L�0�K����7�NX+��OI>`��QuI����_���}G��gϞ%�#�h��`?��C��d	;O�pa��Ʒ��&!��Gx-�YI:k�Y%���j8��w2~WC;�6�>yH,�dti�3A�}q�ͱ��z��L�6���G8��~zn�1�-_˄\��L��c������XG���˲�ӗ�~�{ �/���	�� U���#�-
���܈)L��U�	kN�\G����*���)�ޮƕ_���0���xi��K���B�7�kMoL�i�MW�G��f����h�ꡕA,�u��jc�k�8�x�i��mƄ|ּ����9�����n2G�XSSӷ<��Pp��%
\Bʍ�CMn�8�����q��^�KT��ɴ��!l��
Sީ������y�2�R�����
¯�ѝ�̓wV� ���*������ͮ�i0D>������}�b�LK�Ӿu=X�W�jR�c4�5�MtBC�۵��*�y������������2G��1b*�3�\'� Y+�1�{�&�"��th�(Dw���� ����&	Ʃ��6���b2<��M�«�������� �Ѓ�s������+Aw���,6�B��JK?�*eg��,�X���~��̣��	�7�E8�<yy��i���-'M�`�6B�Og������P�����<k��� �H��sͷ�~���(J4�Nކ�hiɽ=q�m�K�q�E�BM�ݩ�c�=~U�����"�k�k�`�Y�P?|��ѭ#����w�@�O�^o����2*�٣������C�{�mǂ�F�`_C���΅�A�Q�oQ��n|Lr���-=M*)Q�
O��G�͡��S��^ma�N�<��U~-Mie�ز��/��h�*�r�'5Z_>^��J��Z�"�
� �Y՛lKƥq�1䎴:�o�Ru�_8ć��w��}��b����[Y)A�o�c%���z�N�p}M]��";���5�i��1A�$��6ё.���$=���в���S�N����z6�O����@���K۹�?tu]��mV�"���_�� ������6�j�]nĕEv����%ie��8�"��3�k�A�/�xi
+�5��W�=�~�޸�C�Q,C��G�� gY��A r]πN,�{D�)~f���n�ȟ2P[>�	�+b���E��� s�̺)FW���{Ij�~y�g/�g�u��X;p�������z���|Y�cدך�c�R�����]�B��a�������$ء���,����ϝ]
,�Z,q��\q3	z0�x!����7���Z0m��d��n-�F�[��)�9�7�JI�{v�<��C�,P���s�U�6��q�D�w���.O߷�?]�؎�n�����(Q��O����,��	��p,�,_��*Z_c������o������\X�uX����GBG�����5$��`w��U�[Y/d	;K�9�p1ye��DkR��x���-�0��ck�4�?�; n.�A\��[�m����WL��TQ�TI�퍲��lb/(dM�����ҕAn-��d�93����n��*�}��^x���ܻ#瘗x�9�fv�\���	+���9טI������=���D��aYJ�b�B�z��-6�.ԃ>�P$W�b�ʢh	5���$�Fx���,���{��}�T��EF���Њ1�C�1��|���*�7��A�8�61�=�F�]&�]sH����L����U�kfJ=�� dK�s��x����;r>��7-�O�(��H)m�z��c�	Y��7�F.��U��s��yU�P6PH<Ȍ��r0�l�J�� ԛ�i�"��y$y�����Ҳ'Ь�e�y=K��<�;o7g3ؘ�OgGGQMuk{;l3}Ķ��9�k��3�X�-u�=���.��Y5��m�e?�f�,-�+�<�!�k'�&�R-?`7�uR�=��8�xM�g୺���g3��N[��Q._O�@�{�����&���MО[$*��,7�����-�-j�Zxz=>!��bf�M7 �yƠ�� $��'#]�g@�>�*����+ES�QF�Sj�w�	 Ge����"��;��)�ƴ=>Al�êշ,�Y���M�m���C���g�@��h�!�.�#����.w���v?ڌ��N�07ڊ&��48K�<��Џ��H�M�$݀��b�21QQ6~{��'��`E���&���y��J��2�5z��\w�G��_�.Vd��U�?L���Ҟ�<�pδWO%&��SX��~֚���t�B��0<I�~B)BsAĞɁ�������J��g3��U �:��2�ĥ?~���Sa�ɕ�1.01v�	���+�g��Z$�Յ�r&왹8�3���Y�5Rƫ뱧ao6�n���D	И0�E@��:�s�O�˳�������_ ����2k����K1�H��L�B|*�3����MN���)�Z�
�!�On-F���ZV1,Tg
��I�a�*�������g��a�XbCE�Z_��8x���k�}��^!$M=jB��X>�y�;�����c��*Qv»�,�(7܆��r�T���}���2QL�خ���JղC4��L��Օ:@�iBl��ҽ��f�G��n�w'	g��~ ��H�pl�]�>�}ǡ
�7�-,�7c8;����A����"U2����t5G������V֖���QT��g+o��]V�M-�;�ş���`dW��0S�)80�_�B ��Ff`����NW`��{̂R׳�%�QZewz��b�7!z��8X\�O���t�17.�C��/u�����1�u|��8f���}8��f�`�=�p2������2�����e_�m@
�z�K�����2	O���>��R��<�pہ���ivp����ո��O����	��f��Ԙ$(5`�m��v������+��~����F�|u3�����DkRH���Q�����}���g���.v�w��Q'E�0����=WZ�b�ٷ��?�/K@�y�}"���5 I�q��r��G����M[e���܉if�(�S���\(���JuC�o���vr� @GXz�|�Tt½:��mQ�����4ȡl9�~Jе�s8�<����8l��%�ǉ�Yi��.����8����Z@�q��z3�P�������(j��^	B�آ)��\���Yk���j\-��T1��Qz��~f�(p�͎0����}Lj�;K��7ޚi�,�.զ����B�56.*�*P�����'���I�;��m�࿷I�A�qޭV�Jd�����Ώi�Y���a��a�b9�X��X���|NL��D���"�"0�(�Sw��	轑��k;��^r��d����9�����m}�S�Ѝ��N��$i/�]��c��9B?����P���E�k��9�CI��
���
����������hJe\���%p���nd��KV�mf��.�hJI����G��?��(9`l`?4��F�|��s���7���z!Z�	��dC�����jO��!*Pfs�Tmu��z�N����j�����`�������I�3����Y�*Zs��������kI�Vȵj�H<�����=�߳&�V�{��Amhl-D�%a���K�Z����*_��m`����?�Ў��C�{� 6��	�^ha�r\��_�oi��9�ss_��� ]��in�1�*������͜���1�(�þ��`�ֱ%c�APel�;���`��*X�톖\nR�4��B[�~�@>�rK�ݮ?�UY��(�F����E�p1��f�!q^��z]��S�=}�4˧�|��8�2�U��Wvu ���\&4[-��-��3�� �W���V���A��ak�q�?�[-����yo��9�w�X�����3��Z��ʀw�S�}޹�**	�+dC�;|�W2�PhFp�B��b����#>�,�T�>�3mR�.�dզd�'�6�'>���L{�nĴح�2
�Y�&#���NC���:4Ó�<v��&Zyц�L{Kh?��J5�Vw�>?�7�˃��\����ݞ��S�l�컞��!
�ct��^��c4���{�|߾!�
�$e�s�5X�3���k�&6�y/���˘���m����R5��i'�'$�lT}8�s:��Y�JV-��5�-�;'2���텗p��o�"��s�1J�@���E���B���b���.�.��氓�����o�03ޏy�6�p1	T6����""���Z��ݯG�g�졕�e�+�۷%���]:��qSz�K�z)�	�'MhyIN�Cֵ�t*�gk�z������'�����t��s �Z���D+
\�>c�Mb��:t�E���<(�������]�/%J� =��;����/���!Ͼ�c|���]�S���o�ɍQ�?>\���@����a.�K�Կ{}�6td��S�c�w�lWR�}ѐ���5nD��)�n�@f@l��,��Sg��he�4�g��\�ڢ�yC:=m��`�nK��ƺT���!W����l�W�C�Sto��ʚ7�_�2����O��9�E�1�M���������3��٩v;ҩp���Ii�����6�1�{�EwfY���H�� >�u*�}�
[-G�'^�U��R��!v�!�VwW��U��*����51N#�,��G��fP8�XB]��i���ʵ�G��f�����[r��'H�[z,�W ��OT� !I;RE;2�`y��R��XʉG����Y9��ӡk�Pf���܍6J�o�r�JF��8j���o�h�^���W���4�d	�4�����wy���ȱ*=	��'��䋱�6Q$�<"�&ڒ}�V������g�V�G����	fq�x_�ð��
���?_ڹ�o©WoY���q(�z�F��:$�˿���HP��}�Y�����A/g��*�z���4�;��ӭ ����@���i_��Y��NW�,�������<��� �� �^M��+��=y���VW��:�35K��}-�����7��.`ֳo��I��ȧ���:�J�*�R�����Klp���2@�}�
�M�*�ӷ\�.ڛ�>_+�B�9M�mc��aq.�J"u�G}��Q�>��C�9���7�xtn�����:8�_l�A��~û�����
��h�2)���N�x3�p-G�>Yлx�;DF������^{��ǍϮ'Y�ב�N�܌�c�:���^�v~��Dk��E����~��� �;P��7�R������������/r���T��H����R�j�mO�������D�-�[)R���,Zv^�x�� /�1���D����Q_*p�@�2H���ojZ�;�) w��T�{�B ��|}�3�vݮ��	hއ�C���B>�TV����D*��m�p�ҾmP])e�YM_�X�{ǾS�&lU�G��Q==44G�~0���J�p�p�mt*��RJc��Ix~Ơ���8!�O,���4�}��!i���������%Z.�s�o	
T$�8�Y}�P�f���,��!�}�:��<=��~��,bawEnա"-[�U,r���^.)Q/�Z:�����~Pr��tqҝ�g��`2{��}A�e����2;���<�8Ű��}:��g� TD?\��wW�+�U<4� �tR�![�~�ںm�!����8�mی3_���:qsź�ë��no/��[0���=�=o�e1�m��AQ�=^�V���1-�Q�K!���K���{�H=������ U��S
�S�u�����:�Q�xk���_�-c�q�A���G���w9n��$����B+���Г��R���2�t��Յ�4�0c�:�ڲq�p:U S2�t-�L�Ľdm��J��o�,���Nn���T�*9�����P��H��/ɍ)	A���
<0�N�m3����$�k&CR���{~=D0d�?	��׹�nD���8x�wk�;���#8��ͼ�a=�EK����M�
���*�Q�M��ǧ��!�����N!�� �$�����q�:T�V��l�do��%��.'�05o׽߀����w�:�J�l���IS�O�:O�c�:S0S:�Ȇc��s7��G�7�1���	`�Qp�S�r[�U,�B+�K��˅yOCCk��)ਡ�6cz!�+���P��$��H����B�6��^#�:]���a�e�H���R8!���+�0Ǩ�Jϣ���O���En�T�]�t��(��E�Q}K�� �[��z0>N����)6�M�<����1)(0�$(6ՙ�9+�ְ,����-m%�l��ǎ򍙔.�ηS�,�i��4k��[>�w7_3�M����Y^VUv�����ڻ�(SG�튨�xEFI�5����]
Ə�w�;�$��c�>> �,����1��5��偭u�I�O��5�v	��G�ti9����H�:l�X|���(��#>22�Y*�6[��-�7|A������� {�'._5'��˜�|Q!N��W������;�v��҇�=۾�tdE_�0Q��2�-��$Q�u�;^?���ˎ�t�+�3���%j�?����f��4�A��*��#\Ϧ��O�"Ǿw6cN����|�=�;�5�mD�~����=V���_fe���Vͩrַ��6�E����V����w��Ev�u!�X�Ao���[�e<�s�a��^���Q�U��9 %նekJ�{�Np��yU���/^�����5�����Az����'��8mum*�x5ѫw�M햒W*�����qX�r6�����ƫd6�E�r���ES�]��N���2���#)�eU��V�K����~���>iD/H�7bO7˩�3�d0�÷��*�[���˫:��q2�>ì������V���o�������g(E_��d��{�3*YS4�Z�2pp����~�3z6J�8捬�(��N���7�w�ص��$=�uq�Āy9v�����?�!�_Ƽ��gn?y�	�����	����X�Im��,�(of�*E,��eUt��s*4ވ�Y��!�v?���@�C_�V�^����&��H�kM�ŒM���dQI��5���~{^�H�v�T�Z��W�� ����S�i��4����C�e�l�?�������E�g�p�=��v�Tь?j�O��}�Y���9���혛�}�������46���g@\lݭ�*A7�$Eߜ�����lhQ�|�*Ƌi</+��\@�meՄ����0�'_�5��f�xw�xʔ�ix�+
�k}�'v��M�:���;��Q����!��^��2z#+�jP�}"�f�'�H��џ�����-��!�)���t~	@)3L-�F�u@!��87gN�
T��֫��aCϒ�H/�{*qQ#�FNB�#C��K�K�f`�m�'""�e@>�����\>��o�I}e���b�R��J/���O[���8�����A�2�ϟ(Z �l��2+{ȥ&*i.$[t%��f�Z�1,a�!��
��6��+tsA�k{�+�4.Ĥ�ATl���mHC�
(��c@�v�[��I�m�m�6OjͰ��c;@������k0�
q�t󅯫dd��������^��?����$�ɲ�������rV�Nĺ)Ֆla瘟�iCY?O07�&���	nV��%*ձ?���S�90�oyy��N��	$%%��WY)	
��.��҈��$�
NȒ��z�9L�����0� ���D4��<�4���he�o/����n�2ƚ�I��v��.YbR�?t	�M!˃�%s�]^�QE�������Ҍ���a1_��8X��o
bX`by7���|�랫����@��;f�@s$�,���B4)M2 ��u���� �w�w�?G@�i�`�퍈Z2�M�7=�HF�4�f+�����`�;.�0�E
�ū�X�{����nJš9x�%@����.*�sj	�>�*c�B&_L;.Jۉ&\,�.-}���̳��n흖�K�zE�~^]�a�"o�8����;t�}4���F#E�.--!tp��������=�B�#���k�s���<#͸�e�U���������r��?ߔB�X����yzrː�q3ѐ�t)rP�"���@��������F�17�w�)+���l�����G~����S�7t�/>��a||�yz�K�u�^ ����wf�'�,��sL+'��NыyyG��T�Y�h�ҨK�Zv�J������>}�8��G0r�ã�CF������o.䜈0���嵱�#/K��[��@ �1�g��L�Pe���zM̭*4n?����<�*�n��<���B����|C�PSSox���.���]_]�?����@���@}�bn%�%۴}08q�����cD|Ā2�H2���<�0FT�lf6��=�E%'��yqƭ�M�1jb�C!`�}J٪>�6I!sAť!��Q6��j}g Q��Z�S.bJ`�l�/���R���X�\�`����Dt+b(t�����K<_l;C� �G	f~X�|�/���$A����eq�`�w�#}�S��eټ�КA�B�j^�l���L�@��t��))y0�:�'3D��$���;�J˂�!� ��|��7��	�{
�N�碚�IDщL�y|<P�n�ʒ[߶C�Jյ"ئ8�XU��G(E5�Dq�г����P��[#8�k�뫖�A�)ç����{%�w-4���^Hl�[9;a�C8~�����s���n,��&S��$I�K�ym�B�Ř��b��<O4Xf�X)��Lɦ�;N�D��G>�~>]�"���7�����>��t{������;��J����nL|8���uo6��o	�j.���uY���3p��I��Xi-�x�Vh}�y�`t���M[��C�����Z���[��Jg��;(�~������������ϙA��^.�W�Ϣ�ȹe~$��ޅsw�vp�4c��M�d����tδ���ܦ�����]�_��>z��9�39F������"�w�爫r���{#�p,�`����Rk�p�n~��z�UF��Cc̛æ�rlTE��s����;��}O��q�&���+d��2.���A��]���{�vȚ�{}H>�j�-gM��Z=Z�/¸r�������MR�1�*�h�����͛1E��l��{�kuo�i���}P2%y�����1^L��������z|��Z��Gl�ӷ��E�u�Դ�Uj�HKJ}���w�H�1|P�Y�������!!I���ޖ�<��}�3�W����+&�u�}��M�B���6���:����>D@�������Sr�s��|��g~\������|Q�k�妲�ȡ�!th��}�)gJ�!��L�R��x��D1����8��9�(��;-N��P������lf6u��(�ײW�^��>�j�ѱ�?�)K�zm�����WOU<B73�vJ�"Y��E��}���~ǜ�B`�4��j(���7!A��=sX�F�l��w���r�x�rƺ��9������h͆���OG�������A�
#Ua������� ��*<��뚈ߧ��I��eǤ�i�b���@���6H��R�ơx�4|tz�������]���I��D{��_sM�@�J*:�2�M��Ӫ萛�K|s��mݼzyz_�\�P����W)*�y�$�Ҿ}w8�oS�y�������;���3��p�|���r�Z��Xí�P)�����1�AM��ۆbHH�az ��?�����C�|{���E�jxՂ!�pz5+x�^>Se���:��V���IJ���ܝm�l<%9��<F��Ď���4za�L@�W�%����T)�n�j�?3�=F�d2J����g��JQ3���O�&$=Wۯ� ��l��r�#5i���0���`>L��2���i�Zm6Ȟ���?����r;]c���ϽC)fA��/[5rP���f^u���A(�]V�3��$k�M���߱dY��˽�P>{��>A*�Ggg>Cpl3t�z��jz=�/--m1������pR����tNL�a���Mx�|��w�a}ua@��J���gt1V�Ou�sЧ�.p��,���6�-6 �w�+i�zq6Y����@�{���C������>v�z�/{/�^�����[~:^�pa��c!=_b����]��;f|&Y�K��(w�\t�OW���} ײ�A��l�U�w�T����QA��2T��.�K��%�}�2 �@%N�9���k�K:�ݾ#Msf��s���Fڌ'��ݹ����|�س!�?�w��(��	z;�x�����Y���06_��v�cb@B�N ~���Л�GUT�~���w[���!��S�1���=D!�H �MS(0xV��k�|���	˝�tq�b�j)�>�<j��j�P�`1�<�Dy��xX�{
�h��>�<��[%0!:RR�;7n���F;�ޅ���dq�	��j��mG� �������c/tD�˱�Q���r��M���q^�;��M(���`xؿ�|! 3���I�����(�!�c��I�,��`�F��������fT�_��3ǉ!1�|�x�e�w����'���,b�Y2=Y:�(C�Aq�I����(�྘'c����w����e/H�$��`��{B���Mg���Rj�>OXђ0����E�b��'��8K�T�;�{V��x���U����!0�(�7r��i��!���+'|={3�i�i�Q��V��1a.��ϱ��܁V��b�߄���ӥ�C��L�s�,5�>Z�v-�Ǩ6 %�b)��Ĝ���\�� ~\���h;��Œp�ÜG@��Ɂ�K׆t��M}�I��A3������,�-�c��+ |OD,��{������ϲ<�r+M,�r���&Y��87IH o�&�\@/dK����e4�)l�����:Hg}wz�p8����u:��)�u�-^a�۴p��p���=p�T��Q��?}�|�[��UDDC���4Qc%�1N�x	����>_�n}TI�#�|���kc�I	�ߛW��o�!���`g� :ޅ�]����>���N�+��hv�v+�U�0�����.��cJڭ��
�v���<��$nǜ/e�O!/f�t���� Q\�b2����AZ �̟��=Wz�&XP|p�#��^(�h�9��7���Xz���cT�'���(�^O	o�J������E�U>�o�y������T���y �<���y�
�i�2��T/s�X:T��g2�=~ۿ�* ���1���kإk;����7R�{�3�����z6m3J����L
���$Ws�1\fֳ��.�㶃v�t�O6t�XI��dEױ�?��a>�8��G`x]�W�j�_[	z�<(<��0����Ò"N
\��I_2��r�:r��H��S����X����32"��-�}������:t��e�I�V2-�o��*�m5�z�e0ض��_��A��<U��w��)�%���U�_�(�=��̪q�~{1/}9�eII�Xi�]~�	�[ۙ�0���М�ܳ�lũ�fa����+bn�0�%�g�e���[ߞ=9vz���ήM}!Ao���>����Tk[�1�}����B�a��g���K,�\)���f����	�A���I�D�zќȇ�SO���i�c&7�o5ӖhZ�Z�Q�>~��4O%����S$�&R�=/9��2��ߋ�E���gW�H���֔��Gg=��ҫ��[lT3p�ܥbP[��X��:��$d�r�Qo��e�|��c���/�Ҝ����;�p9z�H��}��`1J��vk�qG��>ߘ��1m]�G��sj�<p�N���u[�}��9��Uۼ��H��Z����s�8�����D��������uY�g�v�E)X�9x�/@�ů����7��\E\�ͻΉF{������%Y��sM��D�ѻ7��]�t�V�%N��z��a�l`3���il��!Mx7kV�La�����Y'���'�˧>��ξ���XK�6H8��|���������48c���!#e5�����hY���%d�&��r�'�a����`����|/�����j���|z��S�M�.�
�:�Ay�)*�O}K�}���4ϗ"��.pt��7O7�����tQ�CQ������:�Z�����/]�N���즀�h��`.�`�r��zΏMJ]�T
ڣSL���p�/����֩M�n��0�y|܆�n�{�-�!k^�?,��|}3o)u�`��[�q/zAp�E��|/����i�nx��HyϕU(�ƹX�2����crd��]��q���d����u�h�F��� ��I����X݉7BqTK�����ϨD���NC'��|<�6�7\[��YJ8#M|�������T��J6d$��L\�hO��ҹca��h\|f�{,�Z��[���F�ά�(��_;d�|�y�cu8�Q�n�W�/@Q���#�E�������'�gs�Զ��|$����Rh?�-��b�ai��"���*v��I$�Q��ڗK�o���FY��� �����Y��f�����]i�j��0�ಝ���m"E�I!����Z�i=�{K�bi��4�e�T���6�))�ONp1���H�?R�i���o�(7������C�wD`oH�@q�=Wk�О�|Ǎ�z�1����E�55���Ϲ�o�I�Gi=!F���}B*�E�����O��\�,:�
�M�7F��A�kuzv�|��qke�
��4;h���дS�
�mz׾{ ��P�s�����D��dB>u;�^Y,�'}�jRz����1bD�����+���B�l�.ί��[,1�@�@w"��w��P��=D������;u���oN�M�V�+P:]�	(�'����C��u�q�/i{�1���d��956�3�����"��t:_�L}�ؘ��b1h�
�F���^8E�HLJ�K��&��y��
�����?���Sx�!ђ��IU�~�����S��-�I��ۗ�G�7�ׄ�ƣ�x�?���I��4�ż!�К�z����)�!D�M�}u(Ȯ�C���B�xV}�����-]n?<p�Tq��=C��������B\��	�/@�`0eͷ�6����/]�Zg ��,{�B_��j�?��"������υa-Y�l��GDD��/Ҹ �8�a]��㠁#ѳ�������g`��h��W��Üs�.~ܙ:+H�]������j���M|5qm�k����uc3F��;,+����3س�4�!<7h2uV�՟bA�KIN[�,������ge5�m\���j�>�nz0:m�u�,�x��;<���՗{znw�|�mY���	'&�~:E@�`�|ɍ�"h8�U�(y��q����ׅ������+�4�	\]sMK}(��.e��%^�~�T[�nRII��X@��`��Ċ�QyY+xΓ1�{?�]�m]-�X��k��j�����M"_n?&)�`1�W�l�Z��Fns��/n2��.�#�bb�uB������~�5�T� �Ic�����qqqՏ������?;����̂Pr�pl�s�~�7!�TOU�UJx���S��D�kA���C�݅Jv�Se����k���[Ff(m��7A������D>D͍������1N`�չ�9}�����}e�^Gk?|�~sl>++��}9SR�����Q7��z������)���1VUQ�N��B�M���M1�]�67�L�*��1(�Sd��Ϫ����Hu|����=��c^�oۈ���+'ئ��+�Nw��GآCo��()̾�tO��� ��	Vݵ��&�o7{�c�߲Ɨ�N���臨�\�	>K�|0|v�R��>H��Q���2W9�_�:���8*�gyxL��K{����b(V�2�x�Hs=������p��q��Y_q��M���Wg�#^�w����"Wƪ�|׃�o����ܝQ�x�I���R� �XL�J�M�~����d����s�+qN��J�(S��sc��9�c����$���!�]׸��O����$���ם�s���?D<�m~�1-Z�ߝ�E���ĳ����D�,HՍʑ��Xt�i*�8)�d�H�^r¡`(�9��R�@�㘏c5�S\��VL�8�$~0)=n�;l4�wav�P���d�O�����Ko��%����w�{���#��'�ܦDz%�#��QǝG�*9i�/����9z���U��)wwOF�Q�ƃ6f=>-�yD����q����Pu����D%[�(	��J��*Tӆ$T���A%-Fh�eH��l��2Hƒ}���2�f~�ROO�{�����ǹw�y�s^�r�"�R�(��	i����N?�DO��Q��o�_���諅}�Wl�H:6��S.g�.�;o ��8^�`�	��I>�w9}�k�q���A���s�y�,S)�������7���m�k!�ե�/�[$>�}T=֜)�]"A�'d�X�'�=������b�'y {]���9,���h�X$�0���'cMA�R��ٓiE�7�(-����rS�R.5�Snm���̱㓫��B�N2�йW�����2-%��A��8�\��L<H��S�Z;V�)O!�2��G.������������o���؋�.r��e]�J*�̍�ش�bR`�87>*
z�K�;w�6Ğ]B���9�H�c��p��r[�M���,��Q��ev�晍�}�x#��;h����X}��X�!P�����8	�
 �,��,N	+R�iZ�8�Ο8�xT������fl2$����aï�����׍$����E
��TPM}I�c15!�9��F�^:'NT����#�z�:�0��lE���
�����i�|���h���K��(9��EK�&��L��q���w_s��}2�J�|u���GW�6���Ls
�r�-j�l�u����]��j�=>��G!�S�*��U��Q�_w;<!h.���Z�.����@����w���%d���M7s���6fۆ�93��[�QC�/��fa��>�I3���
AǪ���~�b�`�n*����1���5X�;��l�0�@���s�����/�4M+��9�����`��G�rǟ���� �B\Q�򁓜`��i�j�C4M�O������f����8P<���E" U8)�!>7�l�A&#��R607���P]G��;p`�^�BRIM�C�6�W��:�O���g��ks�w����v�kЩD큄i'a4ݎ|$���a��������@LK�O�AL+� T��^t�/�e������Qsu�r�y����4�B��C����Z�v=q1���χ݈������sk�a���UE���`���$�>���������(��pa�Ip�o��� *T��nw[�AD�ʠ�C�;ߔ[��d݅�������d�:��C�t����3��1��� �zi���&�Z�%gY>@�y�ѩ(�K
���v����%y~yA����pY��]�Su��~��!�`�iT��Az����9�	n@e�)Q�z�&���樦�~޹�jE֌_��N)Y���:_AX�Z��(�'9Д�-^��5�t��q�p�r9�1?n���1�L�ٞ��q�S�|G<�����[��ek���'�<�ʁj9ߒ�_#�g}I��,���ʺ;q����g��I:e��d ��=9B����Fl��/G���Ԋ���j������p�pz *�=@o^|ɎN�DVd	���|����Dm������Di�J�(s�@��Ld_Rz����Vk4s��x�+��~W	N��Tg�����|�l�@A�Ӏ��{�s���x��*Tr�Pu�1̋��/U;A��S���jo �����5~���x⧾�����\7q����x��O��Y�<�=`b�P�/�O./�0w����`t�{�d~Z��5�*#1�x]c�]� ��2M��~���G�{;���Dq?��(e/��}��������?*|3�GT�0�ew��Zi�������e���`�j7������O����`�a�7�)9pv��<Z��<���i9�S�i���҂x� �U�]��z�f� ?D�5<	���L���}�]�5!{�솇lL�����Og+��7$zj̣C1eK�����4�{�^��U�A�-��R�kK+�k���rϽ�����!TYXN0���h�`�-��4�s�-����?OLܙ�_7��z�����H���ӻ���9%����Ԓ]5ks��4�9%�n�d�����2�o�B:���6�Eݾ��$�+w�|�l}��8�aE��d��~�Z�8ܗe'��*�>,�V(%��"7�q�%�"!Y][��|�&��R5+�\U�S����k�4xZq➨ΰ�!d(��/�ȧËki��엞0�6����=@\����Q5r��y�������jn2챂�����'V���qչ��d"�����=�Q*�8����1VNX?y��Dǀ,�"B�*�Z��;1�}�j�ӧRJVu�j�d��6~���2i�Ļ��g��XFу=�#�k�W�4��x�׸�
h�d���[i��)5-!p������F�M�wE~�愾w�ُ
]��$,΢�4Ŕ:SA\��k���^�gD��p+Z����C>��g&jŁ�i^l���}�G�/B�����[Q�����B�+����!�5��F��&�����r���wza��f/��m����.������˧ߌ��@)�����]���G��\�Ou�j�����Ü5�?'����3��LL�b ]��X/�����3$���$,8�y��㻗|Ga����"�l���.��O�&��*[����V�#���XX��>�~ $�����q�����}j��y��o��N}�� �?����G���r���1sv��`����i������t-�=ĳz�u�F�b�+�K�b�guO	�S��v��0��&4�ީ&M8d�mj5�*2eUH�TM�Up��a;���.��6yζ��ri5PHט�Rw=OD���oE�~ڮ,߈�R��6�v�9�~��v5�Aj�<S�š*����ش[N�/���ܝd�ضT����������g���������$��B�Ŭח�m��*�����}�	a�b1�qv�M�n�uR\�e���.g@���R�U<G�y�5jv1	�M�S��|ب��E����S-��ȳڴ�=.(U�7�>��B���b�($���m_������?q�3'G� �
z��&��Ld��U:�6YH��Xv��(1l�Pg�CߥW�G��2o6�k�;�8g�l�'E�S�s���DQə�>���g���o�T3�H3�����6�H���"�OM�q���O����N�������?*!�t���5i���=;���`����r���kb�	�*�H܀�����c���W������7��Zy&J�������r� 8�OBT���8��D���N�f4�ӊ(��=�6���K}��~��S�����:N��d��_�Ui�{�sb;���1��B�y���Hpb���? -�ʏ�%���&`�'NM��]�0رg��E�i��b^Ӄ8�;� ���g(����4^�zP�	�z���a�i>��+��j��L���d�wt:A�?Jok���R�B���wg�H; �5خBf�
��=F!�Fv�"\Z\��߽.�b��2�-��_&|�2!�O�����Y����F<�9I�{u���8�@�"VC�J1[�ˇz/3صvQHW��l�4H��ރX�ܺ1[�ɘ1��m޲��Io���#P.Z��9f�0�lSIĚ��]��F|O�G�I)0���z#��p!��$����'��#��<��-���T���K�`������xY����<�6�8�yzq~�7�
���jf��W�B�C!R������S�B[��2�3�����s���i�5��朴�Y>�C_KC�_1��:�'f8QHbSM�5�]��O
JrΨهѴ�����A{&�\0��#��V�; e%k5p���lZ�PQ�ǘ�����FH���v�������R��O�Wq�Җ����FO-dÑ޳4���/�L��i���m)'D*��\�����(%D�_���gsc���垀^�zjP�����=��yٴ&U��!ϫj�4֧��[:�Hm�vE�q�=��y'��$�����	�%y(��t�7%���c�����fϘ��>Ru�|O���7!;���.Pə��Q���1����fOL>C��øI�� b����LE۩��x�0n'9���Ge���
eG�-�z����G7��=���)I���{�9�QQ���+O۽�*mW�V+Pd�s	@�vՈO|!�'�������ׁ.��w��<]��p�$�N��ܯ�
�쿣�D��_�KU�R��e1����{��Э����w{�����m't�����E�Br0�}��8�=մbnO|�@���Y<���W/�q��~��}������w�+����m!h��?3g���
��({~F�!��G[���ϻ1�J ��h��o|�s��&!�#�
��9Z�ýd)z+��P��,�������K>
�`[ˎ9���/-/����áp��P�[�����7���QV�k�<��(V5W��S�[�IF�(�$f�C����>%�U�җ�H���"��.	9��2ߥb���Rz�m���x��oZM��%!0c�.��|����4��ͤ���N�����T�j��z`�.��	��s��ɏ�K��z��7��gb>-ut:����#Y��5����-�_o1A�R��m����J��1�0���������_��_�y�|����{���Ժ���d_$����҇�t{RW�S�+i4g�*�����xK�B�!�X�%� � k�,�(�Q4z���N�iw�-H@��J�4-�ٓ���A��w�8���[S�>&�:����o�G ��L�CW��v��d�7��A�v�Z��]�:M
,t��U��w�P����K���6ᮐܭ;D�b0co���/)���$ˮ������I��#�j}_��shE���A��L��}�9E�ld�S���i]#sȔ����^�8"��v4����,�����#F���%�]zo�﮿��A1�U׃c-�����ۚk�yn;2'��QanT~�+�r��������J�6�N�V�I	Cx8�J����q)u�x�cH�6ѩh>�z��Fȭ��1��#�e"s&��'c����c'��w�4uVt�'Z΁��3�N,�i�Iq0኿��-,Y�x�+s�*๪�HN7���2�c��%{:j|?�O�XKwh�������q�䜇�H���D��#9��ƭ��<ӯ%և�6%&~���@2֪�f��*�|+�;�
1{&��B,�* �f уf�i�~�Y$ }��p۴�h����@�gW+n��*���ёx8�>kB��<Ō�i5��ަ���O̝���\�c����2t|��5�7� pp�^���
�h�tp�m�H��.���%С^�S4��$���{������x�C_K)�����.�}>�u@���f<�B<�g�*����%��u��ؾd��u#v̂�87� 4$�z-������Q3~�ѿu�NF�.�Y���*k�	��*�n5��GQH5�T�b���q�}"v���%O0�~M^�[Z�qi���_�5;͑���]J���'���L���8�bcp7��sH1��4���צ�@��`["c��^����V�M�-և9f�PTQ4��@�T�LZ���~m=�i���Fy��7}�j�F��A'W�����W����'���H��xN[�*a���%\kl���;�r'"H�UgT����<�	�/�3�F�$VC��c;���
�����W4.��2�!&8�^b�<ϜǱ�GS{�㨙d͇��_�JAfmF�)KE���d�e��o��=��$"]��ӹư!�\+$�	abjnw��2H��jU��Q�Ew{���v��K�r�����=+]��q2�ys�9��1O68�uz&VCF]����禡�e5�him�W[K2ϦM������|�_� �dp�N�Kz�OX�����,��Ko�S}������S�VG��^���7�/܇a��v=���SG�> �(ݙ�`�:1�cv��KʰՅ�n��Bj���3>�������_�7ls���MשM�h����e;�q�C�2�g�>va���}Y�gv��%���2EEk���8�j�����u�EV��tFg�[u���A��y���Sqz\E`�+�j^�"x��eK}�j������������'њ� Y6����w2򊽕��ȳ���J?>�����HN��)o�Ɨ�cmF�f�V���(�;ĉ��d�A8�n���hŰ���]��	�ɇ��S9G&]d�^�"��*���H�+PM1�A���)̀y7�y%�ܝQ(hu|�����F*�F�����DG� ����V1�����y�*��>��^i;d^�y���S��1<���>t�_i�#h;&��CY�ċ�~'�����gT�{�RW�m�]St�?��mxQA+�J�=!G#�u��90��ρ��f+��y�vsBL��Ԙ��i�G��=��j*����?ω���%(\:x�(������-�M�=]u���$�R&�Z�]�]��c!�K�����שD���u��D�U����***����1�݊�-�/�ݨ��� ��
�./���&�y�8A�L��|�L�u{�Ǝ�����q?g���;G��>wEF`�pq�+.|�?�n1v�����\t�Ͳ�*�4������LHH��(��읬,O:X�G ����ÿ�����3��Z9�$�/Xm������~���muQQ��rD��Iӯ}n�z�S�����X4�At�������=8dؒb?S�����Qd��p��в Nmub�qή��E���$�3<�36f�����N�GH��0�^�����;ٮ��AX�w�ݯ�q�N���9�}N��d״�69�D4�gL���H=%�N����C�8�L q$}���5����������\'M����]>�v�"�x?��G׿�+�y��k�=��V�[�h����>�t-������Ih�6�"<Q�\���F:�d�0=pk0 �2���t
g�!u�۝����1��=p@tqv4��Ǐ_�e�|�H_��,��)��������)������X;X6� �WX�S֜�((�p�����
�]ݾ�O!!
����d�V�#L��"a<jFOT%~�4.,£���,r���ԫו�\�b���Xyഃ����E�¯>gס�ۦbjιf�4%�ڳ��|��\iP-�FjV�n��ɉ����{��I4 ��u�/}���aCO4 E�]?{l�H� ��Rrg8����OH�)F�2� ����j�l����h�]#�w��ߺ�RV�[.|� D&�tm�̱��خG/7��?	\@���p[��Qz�ñ�pZ�(�"H�&���/�5腌z�m��_�v;�
�"m����AP*s�9�Fs��~%�⃴��D~��;��h��h9���t���7O�	[Ӆ�]{�r�h0�Ƚ� .�ҧ�'���ÿ�k )�����f:�����'�ک��ls��Cv9mVh�K�g8���4Ŏ���N�޼_�0gl �_-.'�k-֏�^m=_�DUљ�r{!���=��D�y������-IA�V5�V��(���ͺB�]ˠ��m�AHt��o��|�*�B�o�q�)Fs�S���\�a��#����U��^dC�}|�;xT"��7diL0��l�[V_6��_�F5�<0+9�<ߋa�XfC�{��<A���*�:��zߎx$3G�߰� %z����61�m���H��#4�k��Zf����� 0|�?�L��z����	v��z��=� >Z��,Oy����f�h�P�~��ך�GT��L����_r���g�3�ٳ��ɄF�#U�0w�4\	�sk%�b^��j��9���bC�"�����&����c�����C�-v��b?��#o�T���\�}ctKj]�������7��楜�0ȍ�Zn׊_'%ٖ;:.s]ab�?1��^���==7~'����`\*<<�x��.?d�p~�O�9��%�^,��|���t���\}D�x�[�17A<֑�@���l�����+���������փؤD���)T�&m����!j�yهL�<m������Xu]]�(�� U����w"}����mE��KX!�;؜�'�w#f:l�t&Cc�����CO͞�&ܐ�����Z�����F9Cp�u�s���+YN؍�"e���~�m�bZ+yk�ß�$8�Ϻ�O,M��@�(%�	zY(u5�V����Kh�茑]��'���U�.9Fn�i���?���Ȃ˿� '� {���~�0��X��͝�ps��c)�T�ݻ�w�F�����_�a�C' ���H�������� ���$
������iE7A��+�Bn~,��<�{w���7��M�]�8��ʦT��n�����b�밯!�԰�H�-��@;�n��AZ����1d�z�bI'2d�&�ow�h��_�#�o޽ӭ�D�,3N����S�3���s�0���:��O�ߊuƎ��ؑ�AP�������e ���J]I�
$�p�V$%Ih�C�# �l ��0��4���ς G�4ð�S����k=�J"�����9X��Ma�$�m�����`S]�r� �ڱ�#="�Vy'�������C�&��#�N5]*���|n�>������pVf4{�N�m����VT�ȃ�@�j�Weon��B�!�W3g6V��c�������8��*�w���D5�W��g��HM��;5�!2�W���"�^v��'��<�ʎ�}���@�i��i�jm�y�f�y�җ+����b�Zp�pN{��������w��o��yr�������@����tO���6���xŢ��c�fj�
��ڿɗ90`��"5���ަ۲��5��Pg�Ma� �g��懷���ܛg�Rp�־�<�h�m��SP�9��~{܄��#����	Eב��y����>G�»�a�FFn��uZ2>MA��,�D�.,,�?��jG�aL�pK�)���9J/��c[&}�k1��D����Q�l���"�ůI��Ѿ{���K��(����3㝆-�f�9)�,�3�,|~0k|�^xxx���H��<h�#lO�s�F��FA�S��@<�|��OZIIi'�lB�a�`0�b��Ν�FT��H��;O��8 ���c�Y6Mc�Xy
IÍ`p�8����"���� i27F�����|�'���Vv$t#$��k/�k��:S!�6����	%�{�+-))�R��j��|	�ן����Z��_lYfl�h}��>2�BF+(�ӷnݲ.+x�pp�lҰ����U�?�𵃠�H�BI���6b�NE(/��F� �����?֏�ؽ[��˗�&�E��T��<�}�*�c����2�����I"h���&d�l�Dg�U�y����Q�b��D����]�����M��f�㳁M�'�D�\G�ڔ��Be��X��:{��m�Ȃ� ��
p3�z/e\F�S�}ς�?>�.-#&N2�0%���~H��o��?f��e�'i��.P�	����l�rҬ��x/��D|����jۧ������[�K���o������n��Aѕ��+�`6�T��xk�.�/Nˤ��b�>Hj>��Ъ�Q��t0}ͺ�+�p���NF�`;���6ӄ�TC}o�j�mM{�S��خ#��	�d�[lRg�+�[��r��
)��_c&$Jͽ._�A�*�����lBg�}���O,�W���o�8�k��ȳg|i~F�&$�Kb.��s/����B���\�������4��J�/F:�����G�`c|��[�YC��˴`��Z��鍺@;��ȳV4�UOZ�w
�X�΍/��~��k�E�<Ԫ3�\�Y���~0�w%��a�[W�Au�VqK3�>w�M��t:}�q\ ۿU<�ƹ Ε�h��t�L���n��P�g�p��_�s��j �y���c!c_i��r��T������<R���������������@N��`*ԸĮU�MW� ���%�w28�Q��1hb/�; 5Oo˳��zC1G���'�	z��4�[lWc1�u�U1�����R߿�8�-�4�0ʺ�i�Ԛ�`�{�+��b��̿���{��TTA�Q����\�G+<����8"j���ʯ`�� ���9�����p}�^�&0���\|!/jtM��ᱬ�=�-xF�G>�����E%� �+��W�P�@8 �X�TJ������r��>k��5�m� �[�1�� �O ���̷���Y+��b���7��>����NnX�v��i˶�������-�,d�'��YwQ��R�e��)�N3������w ����b|U��- s���?o\:�����V��'s��r��e�u9�zd=�p��fiM�B��/�֢u8%���y�pU���_5��_��� 	}8���6�֙O"�6��{$ X@¡���Q���m�H��y�̃J$Cg3�	�o	^�A�������ÛWK��(T��G���D���Ir��� P���D�;���	`d;�+z�,���G��Yr'S!�?��Z�U��P[	�|��E� Ci��g�)8��ދ����D�/'�����p�HR�0�mJJ��ӧ�V��K�I�vx�������~ҾD󼾾Tss��P�K2��2�?X�~�˦�99�ƹ�#ԫ��{�ua�.�;�j�e�Х4j��D�hxW�GUb����ƞ�ȼ����{S�Q67�c�#��e��+�^�S_4����v�����(�0|r=gw��%��1�T"r��/3�-j�'cjVR�Q���A=n��i��Օ+e���E-��YlS���֔z�}���t��	_ٰ��<�l�<U��&����z$f�ovpՔ�����e�DoI	HG�2�x'D�-`�eZӨ8&u:���vNx}��F�����Y���P�
BX<)XG�9��}�.JER�����<5|mh�.O��aT~�,H�/��x��*���gv5��T7%Y�̼5��$Y!��)���'o�׹�gl�(a�Ay��vBŖ���h��^I:5]l���%}�>�x�̓�G��T�6 ���I�-�n����w��-�.��|葽�r��j��ؼ9�`iY���ܱ�����[�P؄5�G �d�7)�t��܁�xHT��Ҥ�s5��ψ_����(ڠ��"���=��Ի��l�܅���޷�J&��0��G<�����p��;��G�t���>�i�jZ�nRÞw"�߼u�`8�~��k2� q'�~r��Y�2g��z ��f��/�?zb�{{�2����ڹs�ѧ�P<��>p������AW!���R�P�U�w!�w�zCH�����Qh�	���Y�z�>�Q�E]qk�tj�7�n_F2/	�Ϋh\�M��k����+��J������"�-^����+�s����0C��kߝ��0]F���d�n�����䪯A��������O��Ӵ������~����{����z���P���i�5]�}KVD_��tv�D��yeT�sF|]������\��L'�j��ɠ E5|H��n��ڐ@u�P�����70I*��oE���a߭�@���&VA���FR�x�9�U��[�L��m�I����H���C�9���{V[���Qk�"9[�����j�;99��P���$�����=�ƚ-ym�fZ�i�wX)�knL�u��ҝS���2K6&��3ɨ���A9�x�8Y!3�G�#����d�c��m��@�y��{=�)�y�������-O*m�l��z����Q��l|9�Ҙ��ŷa�H�$Q]VR�ō��t9Y3zϻf&)?�Qd*�����䓣p�\�Lm3��
�x1.\�<R�]U�5_�wU�Wfx���
A Q�	4]a�^��Dkjp�/3�p_����WM��D���pj"Z��������W!�8��q)
5" B��R�}�U���k��Uy骿�����r�6�]�I�j�*w����y�W�}Ej���Ua�R>���ٳ��h�Zڧ���:��ؑ�xy�n��vY9���3��`�׎��/�7ФVK͋���XD��_�A��5ر_B����]�/�̪`�0am��3k#٘�5��B����L@��D
�\�:���{��7i/΍�**%��"�kTBqG�v���Q��;$�@�o�v���E��&1SJ����t���t ��Jkg��ר��0��Dxu�L���������/%��C<�x`�G�?}�6K'�3�����FtN�ŷ����oWpƔ{k>�M-���S&����a��և�]y^r�Gw�2��K?o��I!�a�"����Z�,~z��?����D���>�ƽ��]���D�i���I�����+X�Z�P�Ļ��vC�H�j�z����mE��eI<�s���K8�:��m��1�y��>�+6��zT`Jzw���s���[*��|H�*��&��U��q��Jv��V����������C�1�g�t4���m
�`���'�O�<�_J�qs�̱�΢�S�2-*=�|{~g�����z�b�x�~航x^/�<����i4kl�Γ�(�Z9�T�-�Y/wy�a�­5�PP�$��N\C�b�s��_��8x:�x՛�x�4	��$��ӧ]'�Ʃ�M�s/�ٿsxjx���|0�r�.��y��¾7@%��eό�~I�M��4���x�m1�8(��<�{�=�?,+/Ox��ի��7�����8\"��2��g�l�i��"�ӊ���lש��%lD�7�Zn�68�,@��2��k�hFB��Zs���'y��~���w��7 d�>_А��}r4�OV�(�'�d�~R���d}�9~��V���c���|֞�|ㇹ{�r�Q�k���*�}#��N���h~ﹱs�`8etR3��n�J	|�h+l�/:3B�[	4��~T�V�W3��C��N&��"�b�y���{ϔ+ѣ&���6Xt��G��p��yw�QW�j�΃���kK��~�{bZu,���K��7nF������W8�*�9o��}?J��M����ܜ㫤��aVH�$Oc3Ü��I�dN�DK9f>���`���Ӭ��.�qC��h���y>�_&�1�,��B~�������M�9Ѯ�)I�WUA������؈��/_����Hz��H�Ϟlt�0l��XO3���)����ݽH�5��b��zgH�\�m@cǷ�Rf^A����o ��1�
 �$�a�/��"@�n���J1v�me۞*ڌ\��ώD�!� �I��W㊏F_ysHx�+g3�Wԡ.\��b�7�a[�*���D!͊�O��J��F_'aZ�h5,��ئ��o�<�:��'��٘"�T#u�+�w���=�;<:����3CTTT�>��t� �6A���
u����U]tJVF��?��J�2L�J����x3^���zo�C<���0�|�,���룴$w�']�A{l�������D�x4]�RI����A��o<�j�g��X^|������4��	�S␶߯63ޙ�GJ؂;�CAD������7���� Χ=�#�T�������g�o��Di��C�Y	En|۔��fZ�W�ߪ�pi�@��߇����vSsFfo8d2�5e���]���Z�J�c�#1��4�.�:��X��-j6v���XD�Us�3��޸HPX����PAŠx�^��d��*9�C�۸�iӦcQ���v�9^���g�ĝ76�n�Ti�wMv%3޾y�ldd�>5Ӷu/��$\Ck��m�#����(ߋ�
��ʓ�MA�b�����4��[<+�7HP�L-+�`?y�l���kܹ߯қj��}�wE�B�U�^��������G�V��w�����v�(��o`�x7��=ښ�Ig՝)º}$���	�kBEޝXep��'e�#���O��'d#bCC7�N�F��S2����\bl����?G����x�v,!�9�Z��TRO����\���{����+p��۩{=���F�p�;�����2��=4��r�q���ƺ�p�uI�SS�^��KX�/�@n¡]�M�>g\�?�69ٖ���l-e�0MK�����oE6�U�z�}��"��:��X�ij�E��
]��W��gO�uF���v�_,ܙ�8�5�-E��4��y0ͧ�zp��u&�m���u8�N��-��:9����nj�dk}�Q˳�����*0}{�1}��v6y�$T6m�a�OP	����B֩a;�����d�'��?�dpo�[A�4"��"������#<=?/>��R8}��)�bp�#:܌��'-��-���a�Q��F��8Æx���Tأ�gJ fQV�������'z�H|q�6�r��/K�Es/�hч���r�]G����!vH�J�9?�Ǒ'���}�{����\��iR?w!d�����Ya%��k��<ء�l�>o�e}j�*E���{~"θP�d����7iyob+ޑ�p��ҙ��u�s#r<��1�X�o\�FK���L�'�n�.y�-ƏK���({޼��Q�]�>�2l���"��;g���׼�8J/������k�
�&ù!껔g��Ϋ�ۛU1�D[��Wm)!F�H��J�>�,�z�����P1���g��8։���R�nC�*�](��F��:RĘϠ����/v&��m��t�P8[�	Wt�y^�D��EFn��Up�B��ʙ�j����CN�h� D�e7;���`�l�����>'9�\Q�BعS�R��Ұ��������m�e�^�^kU�{�E�t��In��7�R�^7H-�X�Z�����o��j�77-\B RخM�o��7u�=-�|�]�F�q���{�x�2��oߪu��G���,Uΰ���[͖�Nq9�ne^�3���$����n�"{��&{ଌ�pBD�6)np����P�}u�f�%6�Uۅ���+&�7�;pƝI��e��t�>�G n0���mR ������=��ه�^D��33-fk��>M,#�ٱ]�z��
�^
B˹:�O�+e4����|0���VnW�D�C��:ŝk��gl��N��Q07��Y~�YPӥ�
x-���.�D�>O5�W�,��}�L���Gq�O�C��N@���?�WC��Gvp�%G����M�߹o�qi���w���9�)*{���<����w�M��0��ќ�=�7��`E�{o3ڤ�=J	u���M����`8�By��~�r�@��Io��FeF�	�#c%I����^|���]�Zƕi_��zg�p�k�7c�{�N��M�4C���:Hp�Jl�˕�� 5��Ƴ�*��c%�|Vq;�j[��'}V��׻1ʨ��|yP��VZ�⻙]r-��]�2��M.�}v)�M�p��e��}WΐL��k��8)����P�"zGs�����T��{��e�~D���'vP��ղ��8�4Ȍ�z���U���5�c�۵g��W�B�c�*��%���_�N���x4��T
6��M��5�������=� ^BT	��S�Ps-B������NI��hD��J>Z27W{o�̲�����Wo�Z4��Ƴ��=:���ʍ#�C�J�"����hM����d��7$XÙǐ�}��aV�F���X��,n�&ڠ���@}p҅ �tQgS��`��/f�|q���{l�oNB�oB�Wr�~�nc�gE�RQWW�'J�q2��Ċu�{�|��|��Ys~�5G`�#ќ(�h#֟̕���{C|�|h�י�<>t5~I$3����2B$�C�A������7O��Qں�@�;���Z��N���vy|�kE;�1���2�Fq^�Ҋ�]�b
�{�q���/q/v�襅R�L̏E�v�E]�땛�+�h~��D�˟)9��՞ɽ���4��bU�Ç��{E@П�3���6��f��#�E��#������i�1��c�DR�G��%�}���>���.��\Vٛ�4�dR #���[^��?SG{U�-���0���YL�л�\;Ğ�%�^>��4Z��Dm���%%��ط^O�
�{��c�� P����G���ia qI����Y͇k�oT�l�`��@6����;z/�����]�8����6��G��l��TW �Z�Td��C�[WJ/�`�e�?�'n��#q���U�lÿNə��ƘaI%����.�}N�Jŀf�0�,�j���8j����E5�\�
�'�yf`{���4��MG�_@"�~+���Lyvx�|�]��_p�0��l����^���3M[�i
����P�S8��������j����{KCi�BdM[-�MRl=��@��|.R�r�U�����b��'9}f`d�}b%�\%�Ѻ�'�]�U�����O��:�����2�ڣ	~�F9IE%%�G��ß��'��Խ��|9�=^��+�z����-�
B�U�`�}��|�r`Ɏ���P?������W��]	�6�醈���+ƨ8�$�y��I�j��h�8��N�5�d<?qٍ��۷�:ٸ��3^%�BU����"!��|�d�vJQ�f��O��+��B���uH��8�s��s��`*�(����ʾ+���v�~�~=�ߜR8o2|�̾ؒ��w���x����>2�@�<q�Jn��p���2���B����x"�O��
��8�<N��9��]�T0�mlj0c͚d|�kN%Lx��w�Y�]��E�J�Cj�Z���7!v��� �d��z����5�	ԯ~�i�������y�9t��y���k��]~Er��YK1�e,3w�Y�T066ݥ�f$����O,��hZ)���67�T�������Z-*�v�ᾳ��$�{.g�|&g,�Дx:�����7o��(�WV}��!��ɨ�d"4�.>_�i'��,�]&b�n ��?�7�Yd���Z����e���p޴'�$¨��i�ǔn{�<n��%`i��=7h���w���B�ٝf��7ҩ~��
��aJ!dz�ۚ-��m��֛��X��KXJʞ�ܕ�p����#�QW�d9���
.��#5���j�ټ:2G֑�wD:T��^֗2��Y݄^w/W��-I�	�j�H
�BsHѺq� ��]�5-�m(��))�m���f�����
�"_r��]��N9�8���sPZ�q__Z�vZ���Q�r�0�kNt|u���b)|E��>$�9���s%QMg>^�'��=�-��S��I=�08�>m���
�pB�c�"���nZ6��F.|U��IJCϗ��-V쟝��ibF�D�#pxN���c��$H<�a�5_N�ǵ��G��7���=V��#^׹Q����[��+7���u�Ժaf����#VP�d_Z <a�Gj{��q�������'��I��V�/������ C+A��Ḯ�q�K�Q{���32|3dٽ[#��^
3�°�w���������wB���₵3�G��.uu�mI�{T��99¸V.U�Ec���$.mIY��l��Cż[5k[{�P��a�c�acrV[y�9���JT���>��777?7	�$[��䕕+�}���� i�{.uHs>[EE(�o-�6���\lF\�	��T�i����V��m�NDpf�����S���)����0
_�h�5,�8�4$�ZҞn3'T�a4E�Q�� ~�4�ǟϯliF��I|K ���2l�n��r�,Yŷ"pS�g[��^q�ɟ�"V�f''X�]���@{���e�|��l��Yڎ}�]��?��;��l��#MT@:�  "]�DE�� �*RC��JU�Ԡ���A@z�-�NBM ��Fg�Ͻ��y|I��k�_Y{�Ms��%�to&p�  �Q�?U�K�ו���-�0��$n�w,|�Gި^z_�O�֌g3�c���lc7$(��������6,�$��������j�
n���4��M����,|�ڞ��:u�t�~�!Y��A�"P�P�C�!
 �GZZ�h�o���f�x\g5Ϩk�8���L��}�ܕ������ɓ��
��;zz�޾��(z�!�_�u������!hP���>[Wc
�.dhxͺ-�
b�=�l��Ө=h�w���+}}�=�LF�5�X�xb`{}���xl����f7��P��йR�����3����>���z������p1X8%�5�O�i��g��sM���$��~�j���=|}�Ey��Q3ް��t}1|·)�N��n�<\�If�|ôN���:Bx�,�+Ϩ�
?g9q�W�\��z���+û���M��t J�NP��&�n3a~�7�A;���s�^G}���I�n{Fo�������-���<
���{�������6���\L��x�Pj9]����O\�z�p]o�#���v4��E|���>�]�7�ɨ?1K�e��0�*�8�CȦ�V!_Om�����_��Ѵ�Ut\i����>c)��|�g�G���W�����>9��*�U�GE��5�i�3:�xT
8r�q�+.�kv $��h�\��"�aw��X�x%"�1G>!�]ؓ>y�s�܏>���M���8'�)���T9���UZ��Ô*/��w_�n��%�tI³pu,��s����|�tީ�5 �0�ӡlM�s�F1��fߞ�� ۻO�J�����7�#rS�cSw_�!����N'fsE}�0�N�n�Z��P;!)��8�:�FN�הxٽ<�-!t��]gnW��!i�I��}>�����}��$��d����ʒ�`J5$%[P,���I�[�v�����}����޳\�,�.�0�z��\剿1����C�����O1���-��5;�Fn%¦Uч�S	z��qfPܡ"��3���F�y9�G&am$���mV�|�m��6r]�l�����\�b��!�9�������̇wO�N*�9_\%���*d}�K�����$2C%*>��iΨԶ����(٭������6f�C��s�b�G��1���4��<���
WO����~΁l'�t�N�F�-~K�G�޲:�KA%�����RL��u]� �,sݢ��*t���F�jPd��v)	'� ��s����T?>gf���R_
y��P���cU�,r��L�Y]60C\|�,ę��N;�����O��4�c�}$�H�+x��h@�Z,�k�l���U�bY?��7s���S3	|�^	���ɴ+�K<�^MG����-�t)gA�����s�R�ܘj�H�R#~ɒ?��@�s�ï�CZ���i���t����)#COiUh�F���p����@qK^�;���:#��M��D�G�oO8&?�µ˔-���O��P	��}��;�c�I�c���BUCF�A����W��dQr��\��z"dR�'ľ�&��!������D�y�yj��(i+Z���@P�C�Ů3ߴ��UԊ���=��/+���G����CyG���[O_��ы��qzV! ��):d���yH��R~�2�ϴyC��&
g��C�w����x���q躠�`^BAR�潒�;��%�P(g��`C	"4):8�G!?K���cc8'�?�=7��~��^��(/���>�=I`|��<�T_���`�^o׏���
�WI�Y6$]��F����a.)&Vj�C�ڙF5�c7]��<�c��T���u�:?�K�O}Iװ3�UWǟbѻ_
�!�g�;�t.���d1K����ɒ� �� ������n3����6ښ��xlu�\�B��!P�?�AD�D������n�>嗠�r�\��������WH�G�NI���
�'V�i�I��F��t���לP��i��_>J���g��'˓�OP�������+�=V7�e7�����e���@��-'�}d��= �V
`��Q�;T���)��˷��f`�y�����V�7�D<i�h�qyRE�Ud�~��'69*P�{/�Y���!I��vuc�G�M/2+�<|��-Hm#�	!�����������Y��\�����3�(���ߊ���.C��c	�i�e�J�v��C��#M?嘾�� �<��z�i�3�Se��u �z�Ǽ�3�H>�>��̯��[B����%o��x1�/�gH�Ѩ�h��(���Z�'�\[XLE�6���]���_��]�BI�s���b ��@~�C�o�S��X;���&�܁�����Ll
+�σI��f. �j~��k��ҝ��	d��>ᢑĘ��7]i� �OO1���ȼ���s�f'ţ�49�x;��j�5�P��!		�c��e<Id���4�
����>ؙ�Y�m���L��mO���#�E�)�(M��v2�^� bb�`H��'��kB�-�6Zu#��ۭ[�F}!�oٌ�vyii���/��zGs�f��@���	�@���l������C��V�����#���ӥf5^���nW����b+��&���e�ݗ&��z�t��gNw۹��}��o�rk�I�Z�;��#CEɯ�nl�'�kk�8݃�]t��wU��w܋�&coI䢽���1��V�9Ze�M��=�5��z�z��I@WUJ�H&��0��'�X���ӣ)��� �Q������k�qs����&ȶO+��B �J�򽀸������ ��������o�~�,��u��(=�4���h�)���M�U����d���IF]����Ȁ�4 ����'�LY�]}|rk����d�!�A+l���3ͺ�[���|�r�D��ʹ��r�X��۞�?�� 5�p�ҷ �0H�ډ~�D�r��������fy'��W9Ϡ0mANs��Wn;�A}��������I4r�}[�1��5�eL�0�`o������wR�gR4�tp�r�<�Y�� �{>�=�4K�㖐�E�$q��.�䵽pL��DZcB}^2��r�_t^�6��
��"C���D<
�� �|-���a��Q�M�� �n�H@&��[{�d��?�@�<�|��p����y@�j��<�^=DмU.���������(��m+9��K^R��H'�s$J�Q��/�� �B�Ul
 es�xO�_�Rw5�d�p��B�	��_�J�F�Ʉ�q�fA���jNv� �B�.K��w�<�Ϩ��U5G<>����+��m����" wM�i>& �e�=��ᇛ��u�9��,��J�7�A��eܧ bey�O���ݗ.�6s77��*�ջ��3q%)+�}�aw7�z}�"��9�Ol�7��C�<b����t*��@��ނӟ��M�ޤ�O�,Fl�a���O�ܣ^�R�.n���6��3��X�UH�*L�j������*FN�P����`f�9w�_����l�2t�E�$�f9J35R_1]uSx�#���8Ey܁�L1ں�|�k�a�n+�7%�
���F��'��,�K���P��<֑��-@ȱݔu��<^�tQ��w�Qn���1���VxԈ���"�&�G��\H}�E:4)�IDWu�����vw��_c?��$݉Ɵ*��V ���x��#�C�l��u���������on`t�y��D��;���cP�1�Nc#X��-��j��x�����S wd�ɾ/3;�|#��(���j E�&�0���K�02k]��4�¢��)���%�2ȶ�YȔkMD�mO��nE֭�r����w���p�$��I� e����[�R�_�*x��'��l�Z����:�#�5�9��������q? �6[뛴�$wg�u	��AK��<YLx��g(;`�WҸ!���Q�Y�0.������D��rzy��T��\7=Ww-�A�K?V�0ۏV��<Z��L����9:^������d�[��ք�
�j8�+h@͂'&J�⬳5a��0�+���+�d�7����I���a�,��V��T�}�nb(W:���_�|ч����ro�����1g�I��$5�௃������6�Cc'��iTF�iPk)��>9��pޚL�b�-@?'�L5��9�iHGſ�0(�;��b\��'���=r�< �G���� ����S�|t������)�ٸf�Έ�G��2�PU��������儤U@�X�C^}9MXmq��h��w������Z�V�OHх�h����������P�1��k=�@P Hc[�I�m;I�]�~?�z��N�4�N�uQ8��/��.�\�o/
}MQ�2聁,<p|0�{��a̔�Or6��p�/���&�T���~̋^b�Ho��ħ�Ƿ2��T'�4� �FI�+�b�F��_���ѻ��3��\R���>E���'�yn����^4j�ɲ��k���*���e�5���H6r;U���Й�=����� ��%+���.��R�|!~��+u���^~���q |��5�	؟To�n�O�+����@�݀Fɬf�a{YZ`V���G���7E��"6:�� Գ���n�"�om���	$H��ɛ6�
�S�>m!"auT`��������=Y���y2�U��Ǵ��e6��ڵFk}=z��@�[S��*�p	��t�%�o*�7Q�[N9�x�h�,0L�����d�W��E��|�r�Ԟ�.p��p�obz��p�@�o�&@ZA�Ǫ]b9�ʀ"� ��M�ɺ�}(784�c��!^�j�J��kg��Z��Ϲ��)���j���@�A�9�/<�7<6�g��燨C-���Wɚ�J��p)�$��񝂅���$	�q3�`'�ܔ=�W�?
y��Q���Γ�.a�s��0&N9��w^]Y���4� ����h)FӱWGX͎͠i9���L��A�*�q��+\���v.$%"P�?�F<��FA�ȍ�����>P�D�[�s���A��ϓ
6r�N��ｓ䙫���;9�!�^-�G��e��GK���Ec9�Q�9��}?B���O���m�L�=�B��NT��hxpgy���3��u���X��R4��� 1�MW���K!����tNU�p�����yE�4~��w�Rn#L��nH
X9�f�'�WR�ş�V�gVv1�I��Fn������/��VS�D̦�$�����$�x&3/��x��lh�/�}�C�_2{�2�"��^?���D�6>+U�6Y��V��A(v�����D���x���*�P�6U��U@ �e� �X(춧�.j��f�/��\c4җx{Y�{�cs ��f5�l�	F���ܪC�k�pf�r95��<�E�SB4�AGX�0*�.��g�$d���A'G:�I!�/Q8'�ԍ&���*���B?�3A�����Z��^<SI��FCg�/x�.P�z,�	�܁��}ݤ�*蔵�a�$@Ɯ#	����)�5��/����t�V�`�5���ȶ�ĵ���T.��Dyȷ.�U"|c�k��E||rF��d��pӼmO�����D��2�f`�@��\U��5�Rg�Ws=X��(}ӎN��}S�����p�֨���"���͝3���і��CW��Q���o_��b�� � dӺ���l����PW< 勝{࠻Nl���}�d������V�*��+@�Ю(�b�g���,�K233g�v17>0A���Y7�@?���ᥩO���#a����c__-�+�M��FH��iY���Bk�2{4h�[L[�~�4 Q���8����W�D��NO�T{�����ܿ���z��`�������;�v�oN� �Z�����̸����l-q�H�I�H�Y��V���cN8����r��S�ayI&�cB#U�'`rߣ��F@#dh<H)����� k���NxR���g@�\@�C�,��HJ���"(�.���}m�[��E�o���Oz�[��+������K2�}�]O�\�W"Z�>y�g����'�U�tV�W��ݿ7R������\MX;��#���j�+ڡ" �>�s��-������D�X�/͊�g��J��+�Th�G�z]��d�*���x�x<k�z ��D=ʿ�J��#X]��	2eL_��-X�=����	Jc��+g�x�R�2N�8-'�f��v���G��Ԏ�M�?7�'�N��PvJ������sW��km������*��-�7� ��k�t��J����{��I��/N �_%b#�1<[:d�޴�6�E��ƨBWoj������S��'�2�Y.���`@���ο&r�@�O��G��%j{i�Y���t��S�f��u���$�$� 6�����٭���/H$~.��[��>�����"�����h�8�3@V��M�+4�	IA�F\guQ)�`��P�!�T9X�]ʓzYw����;:��/��I�c��e*��.K#�	D�s���Qi߸��\���zb��b�@�5���/a�W:q�$t�ۊ��8�����F�a��K��MŊ|/��)�z�J�UZ.�;(�r�'�SI���ϭ	�%�6��ӡ�&���7�u �����������	&��	�?��	��O��u�{���V���o�ͭ₶:�W�쉼���e��հU~m mx#�c�ھ1��\��A�(���[ˁ�����h�D�T��<BO�dL4���m��T�=�p#�U~���#b`�y/�W�#Rh�sD���+�����b��:��"�ZE%j��@V�EA�N�5"f0��ZH�3\�P���>�'l�l[�1�ŏ{u�~`�A��Nh��|s%���s�Y]��Gu&�n��[�~�r�|�W��΄���'����jE����AP�D��wH�s�������]��{��E�_�Wܾ5C*��I�b!�r�~��Yp��4���ο:��BTL`7D�����v�eR,��O ��ǿ��f�Y$���T1�D�����n��L��< �v��œЀD����Z	Ta����*��	��h�����������1�UM���j~ug<!�L��ouο��k;ʉ#��#���s�8��&\�d���-�G�_�yI�����O�����_�,��츦q���[����Y�J���3�\�o��C���f��e9�Gv�
n���X`Q��aq�/�l[.�}(�0�3B�U*[+���;�E��o�)����2cg��K)��o,6ڥ�=�_%���y��-#��-���@i�J�5��4��ϼ�|��7d�����ma4��}ro�$�����?U�-ʊm���3\��R(��m�)�U0W�ӥ�����t-��"�M�l�\VD����လ��׸�k4�"6�
�}�����s]�kɴc�~�eӋ�r22�q�:m�P�Ks��[k?1b��s�����ۺ?譤�2&������\yXN�ͪ���U=G[�����F=�νR#W˞ig/1��T4����wI�@���X!�x��	��re�O8�p;�Mb�wG�3)9`wX��҇�!�Z�#m=���jP;t�a��N���Uɧ$��g!��g�<f�[���ï��e[���苪3��~�bw)�E��r���#�5F����or��w�F�I�4�M¤�_���������=�#��K<V�ڱ)e�.�
��O�N�G�TԱUK�� ����5�.�2��O�Rk�M+��x쾦�%գ~%��E|l�R%K{d	��W7�M���=�w^�d�^����Y�E؆r�2��t���|�J|����>aX0'l����.���Xe����N���GƗ�\(�O�Mj(6l�%��;�~z5���eP���i�����~Nw]��� �d���ێ��O�m��^e�!���h�ǽlC�\u��}����T��/�k�]�������sc��N����A�
a��Mx���u{$A�n}�,2*sЙj斑�_
�?�Q�t�\�1�麐�P�06���w���,�I�o�j.>�F�����}��˽(�|M����Ό�6��z����P��Y�D��S���_��]����q��V�c�7bv��`�$I+�l���d)��E�g�l���l�m�h� ���ɲ�"���?>.�iT�3����Ooxak��F7'��s��� 轢�*��'XU����!U*r<l=�<��˴z)׉�o;LKe�?:��|��-�����L����r�H1z�؛
�����{t_�F9�̎^Po���7����C]�c�L�/�ޢov��|��!�K�C	�wM嗠� �B��Y����bi�c���5(0%XJ��w*�13�����^�ŀ��0��_1x�l�P���½��y�b���YFx��鯻 -��H�I,���}�M'��o\���m��%�9x�ȭ*:�#M�C�i�5���g0:$�<'џ:l�#&��Y؆����rW��W%��e�ɓ�d����Nq�j�Ά�P����l�NL�ꟴpg�5��{�����w�^n$��e��>H�c�������>���z��0j�z6��TV��~v9���?wb1�1�bo���vW����[�(�b�9����5����9���b���?c5a�@��"\=��*�@��[#��/��d�6��nы��d��K�~�*������b���z_���-�)��"��/�@�ͷ�eaؒ1��l��;g�% �=���+�✼�Uk1M誔5�����J�gpo�\����l�*Ÿ'��jx�x�~N�-v/�]��ݠ���Q1PF��T��[�i��*�ڷ���uU7��M���&r�i.>����{�(���D{h�<`�T+���D�^w)�<��2�b��w��1�N�fe��C7S�Mnu�M(���7��5o�K�Ժ�ǉK#}���#��M(G�q��2���$�����Uȫ^�oEĤk'&nu���7���~XՕ��ۚ�"�40�l���jA��	�㋕\;��,��wR��4�_?+��9A��kpbv�2��p^>�~���盐+�S���.�>9-�Zz�9�ng���x���so��(�s0'�0Dch�ʁ������N-%i�$��+a�@�|#�ks$׮����Y
;¦�*4(�^����*c����&h��ikS2A�Zڕ �P�\�u�q�U��Tjͧ��F���p/�N�v�	jU��k����B����C?�	?/yQ@%�M�_�'�g�=|�/%
x�����o֡���E���z��x��iט���]��b���;�bͿ��RQ��Xo���¶�5����]?�V$����('�/Ʈ�L��4���~�����8k���1}J��c�I�Ƀ�(T��14��(S,s�%@n�U�xjm������d1�7"F�Y��o5Qr�$�#"G"[�	"+�8���V��iuH�^�BU
�����]Q?U*J*�H��H����l
S�;��&�V���%KC��%m�+�}��3I7G�iQ��̿s��2b�X�Bpu`лv��<{�x���<�j]j���j�yU?'�	�S��ne ���ܜ`�R¤�=�o!TB!0פ�o�$���kYd��|�F��*�~ � �Ll�N�ѳ�\�L0^�x���M��'��	?Hf���a���䅬#��X��� d�̻GCir��f��m�
��L��X��h�kj����ݱ�(����B=k]\�����hW�]IW9�����91�[�]0�Xs���;P������,�1��*����������'%X��#�0_��dw�Yh���׉~)�΅�S��/0WVG�:x4p�z���.̮���ֱϥ?�� �;�G�.c�;a2$���Nv�DJ��eD�._�<t�El�=�;�����$��#J�G~/���@��em�?Z��R���Ǆb��7�K	Ő�q��ei�f%�v��=����-VoO9$3[�C��`��Öp!�}7̿}�y��ׯ���9.eu���f�'�*߇�S�P<���6�V����<��Thڈ��]H���;��X��J����^���>I��ɲ�Ne��>b3�:g��srdl�@��@�@��@���E�=�vg��N��&������>�5���K{�\20�kK�5�����9�r7/�&��8���}�S��Zay;i����P,���AN|��[ JZ�N%*Ҋ��~b�5��8��D�����-��&�K�t؅CLRvf�L7��Ok��ظ'�3$@I���Cy(����A�,͘��`��0W��R�]��S�qus'�Rj9)T������Lsj�o__0e�*'&_�,�oƧ�-���Q�p��s��Uŝ�g徭���@��>�;���z%K�Qm5������!��7�>_����^ߩh�+ҫ���$�#��w�4a��3�g�/f��T����ϙ��@�o�;^�pn؞�|���G�C9(�����pcZ'$r�S�����MV��w;���>���},�F��T0�f���Y>6�*�B�o���{��!�'L�F'S����	
t�<�ҟ���fހLlGt���lE��@8�µ��]�3��c�� CO�.�N�Q�cT�%��g�h�E]�2��Л�Sz���M�쌋�|�}���z��3.���8q��RQ\��b�ӹ ����\Y5K���0� U��Gh��sm��+�rO�;�����5+H� CY��S��}���~
>s�?D�'D�`��a����O�J�*	�-��T�镀y��i��ۗ$	UND��;��ʽU����a��$)�^6	G�R)������)�D��="ڽ�y��Q_�'?�Y?�sj��;��lۜm�/� ��$GF]��4:�7G��h�m>���tʝ�sv�ً�qG؜�5�#}�x����U*�� ɿ��%3���HE�"ym�f�.�c�"w��Xg�[V����μ�C;ɣ��u��� }0��|V���@��Q�?�S.�Ύ}�^�6�;88(޿���f[�wX"�e�}���,| !;�z��	������"�<ۭ_`�ғ��Y]�~���, �������2���O���H�J�6�+������|��i>o�+C@�jd�τ��cs�VT�n�~�j�<&�,Nc�U� ��y�;\�Ȭ�=�s{2n�g1��S��~��X�K^���У-̽�d�Pz㳑��&���� "�=�(��PY�F�P�3}~�cb{�Y�	���"�w$��NSf���0�Dn�-�����س� �m˸+�?��Ky�F�Ps�_�}x�'-�ol
�'�ƭ����P�-��KJ?W�t�s�Ε-�f�9D?��{~q��	Ք}�}������\�d�ؑg����ͤ���\��E��sQ/@�;�����
�'��q��c��`e��4�0k��nn�׻��h��HN�6Ǒ�Le���#*t���/b�m�eέqeӭ�`�Z+}��-��X\��� >ͧP�,e�m��8�TEI��e�f��j_�����]�cY�� ��;����ur���3J*�E�n����k>��` &�w �Ċ\-�㲻��/�Q
1�(������DƖ���C'G�_�Н�;B@e(�/��e����͢�_�H�0EdFk5l�U�	�Q7oS:��a���D��PvB��l _��{�ni|��Ȍ�8z+������v��?%�����"��i�A�m���[��������v��u�%��E��鬻���5�~o��K���	�s����`_�R�	�		�y�@0�l�wU��m�v�B�3�
����yyE@+hD��B;M텁��=_ov����C�οb?9�LLP��u��ו�^��ܴ������2k�C��پ��=Jl��ޯ�3W����rs�
g���T?x�9
�W�t�9���b�1�K1����fY�2u�@���:���î�N��.��6�#l2|V��i�O���$�d�\�9*Q�ݢ������a��ϥk��&X%2Z>�C�K|�@_3^��e����_�~�ld��L����~��7=�P�ȃ^�9�[h�|(-q@xt�D�����n�F�2��q%R?H��|Ԥ����TyZN�a=���@�$�C훝w�,�quz��%{�NO�����3�T���(i=k� �:,Վ���=�:Z֥�ݦ��?�]6�4���Zu�	��w�R�|�~�I�5�w�O��F]�iq�f�`�n�{�N�e���:#�E�:�w�g˯���xnƟT��Y��Fp�K��ܜ�;��n�jPX$�� ۞(��E�8�������i��A��sA���G.t?r{�`P6w�����]	Mc|-��q��E�����g1�6��yr*5�-1��w��f?�(�(��D�sC�>f�+�
}�ﭛ7%S�&��
�m�j켪	ڈ���smT�7�y��t>�l�+P[<ݤ�����r�(d����U��/Z;[��� �������f�Koc�7j��C�P�݇�L�������]k�ͪ�s��v������?�����*�J�Y�(�gk�����Q�n|�1���AM-l��_����f(� gV��xu��>�6=`߫'�PОFG$!��%��N�X������Y9�@l�s��Nh�ݾ*�T�h�k�K|q���Y��_���8~���
kpxR��B�m������3��F��ݰSfC�]!���|�
R;wAx��_�>��6G;7�lh�n<�	�ʒh�-��g�����X�n���m�=?��ӂU<^[����#3IrN�1������.�ڡ(�~���_)�E�e5��dTO�Ҟ�＞�9�^�ԅ�M�5���Jij�\ṩpz���is�]<DG��>9B��4�{�e�mysD^G������y�[uq�+���*�N��`ܓl/a�pC��ևg8I���R�iX��@���� O5��,HP�$|#ٛ�"���b0��ZLP���� �.�QI���N��0��NRmzO������$�R����ɓ�*��G/N:ZY.5�+m-R-r�!������ڹ��-!t��I⏯�������T�:e��r��^�VSDk��x˼ts�a���Ĵ8�]�K	�M�*�P��P�C��΀��-��d���M��$N/d�;�=�M��յ�S?uv��tp�P��t�_G��~�v���m!�ak�^�����+�v��t�L.
˭�Nܮ�'��?XF�-�\�,DxKd3��/{Яt�ǆT��B�Eט!��@��^k?Ώ���9@�����Z`�}6ܭ�&�����p����:��A	��;U�7u,�}@��p�����
c�(ڂ���	��-NO�-�eMj}D<H�A2R-m��.��YA������u/��o���9�N_��%0��0�:�W��k�V�M_�i�Ћ�^PGq����e�~�r%�g*+�Đ ����>�4��!Uz��3��8���� �Chm���hdndn'ܜgaL�?�d���J�刺��J(� cR�����,s��nު�H�V)F�aM��&��m2e̬��O�-�2㷙�xs9+��j�
�o`7*�U��!O�+s���=���9�>bq#̼�W���8�@]\+�KtV�h�{8/��ǔS8E�gms�zi8������t�-Ѥ��(�{�Ye�& �-��2A��ث>H���sD���1���3oEWi�1b�E7HȨB��}�lx?_��WpPl���Z�z���Us�*�,��r�,�[7}���hp,�5��
D#q�/Fr}9^�>0*�b��#�)��[UKٔ���Ybں�2������+��Wg�D�Q&���n���{	�P�����+:ϣ\$dRQԕ �f���,$���3]fk�Pi~7mG��4H)Kv��m�YF�=��SS9��|���̳$LQ�RŠf$�#i3q�q��'��N��E�l�(;і��|�^h��\ǟ�4s���J9�<��f7c��( Ҙ�L���
����[��� ��=?� U�=�]oGv�DqC*<�QBXJ��uu�ce��sA�č�#\�=$V�����*�G��%�� �ι<_G�"��%kmn/>I�������������.����Q��v��RS��X�ty���sN!|�w�b�z���Bjہm1���ZA�&y���e7��e�X6j�8L�}��l��m�7��&��%���ͥ �Y���{�,Km��-f�`��Xy������Vn����lx���9�7�2.�<"(5E��N��e�#G���T��::��� EP�����Nk��u�c9y�J�z��*M�_'�(8Q[�t��6�7
1Zr��v~�Ѕ9�L�߭q��<eKW���p���0�m�����qvHz�R�./�yR���9���&2����mln��6����N�sx��2��j\�#����V�8㻚�y����E�g�V?�YƮ �K��^� ev�%���/"��c�IR�f�HC8���j���`��U�8�_����z���v�0�f�y9����CQ�$/�!�R���� ���7��b��C5���:�=�"���ͺR>2��$�s	��V�t|�~�-��WN)������#�OW�Gphk�d�u�1rٰ������A�z�S�*�Z����Eoh��y5���*Z���Ї�|���N1``�g�9��1��L]��r���N�C/F%��>9�Ŗ�l�W���y�=* ����H����{I�O$�$#1��_
�{�L�q�e�����L�% r�rt.�@*#=7�B3�J�>���"�s��Dϸ��Q_I]���.<��L�����ܠ���-�j��m�E+)���BWzS�|� ��媒M�%q錸�`X_����ː{Լ��J/�D�m�gaPJ[�|�4{��nnr[��'�*B������b��GF(�oc<vբ���J��ͧ
�~��|����}�Ev ��bC����¯e�����:Yw��X���F.D����(^�a���Pًi=����W^%���`'��˾���>_/��	����"�l��%y�k��k��*ߐOr��|i���ׇJތ�8�Uz�N�eX�I��
��P���LO�z-���ZQ:U0(AF��'�6�`���z��o��\FE�Hb&�^\H���U'�b}ߟk7Ql�~�>�X	�������W�<}⵷�n��z%pz���}�$�EkN�ߚ���>|rf16uDsX��f~�Aΰԥ�b���7�����+
܈gw7z�PaG��Q/ة|S7�+}�֊� E)�"�ĥ�>���>~w�HW�8���<���؀(�(���ĳ J!"���lm>��.��K�~�d^����}F,(qE.�B𾥎���j�s|��Z_I��s/���YL�U�0{uH��a;@J%�aY��$��+#% �:%���(�7*��%q��8�*���#v� �S�]S�-gv��d�xw(�7vۆ	0=�?	H`�)��'m]%>�e���IRg�f�W���w4�)!�8l����~)[�0�t+���}PC���h4��s�=H�]�u#�۲�xTT�����!�;��*��=��/v�64pՊ�H�oX�<����y�:}�＄~*����,.����#$_�P��[]��74x�e������ޡ��p�Pr�͂�����5����C��I�Q̇E%��0�AY��yz��i�)��+݇c}� �T��k}�j�	��_N�(ٙ�)5q��W]`Tꔜå��?��p��x��axB�q�m����eevE�cJ�~z݉k4�f1�,R���MZ�����`�|��	��\�0�s>��}�cx�u�%�����aaz���W�����t?(�"��e��J��N�s��}В!b� +�-�=�t�ЏU����R�֙��'�ݱ��G�z��{��]���TF�>fV�N�����i���'��&H|$�%'n���K�7�+V��k��AKJJb�>`��K��*)SyZ���5D�/jpK|�o����?ww�������FT���k����%�g��[�Ж�0�i
�>��m���q��3%VF��H:��ݥRW��ntQ&\$��20�����>��L}X�@��8s��E�۬����Tj�,�ድT�8��pĠS�xo�(Ҳ�B�-5fM�줝������0��{�;}�k����Q�>�6�D�4y(�A�����cz�������N-j�?#�L����"�)/�;�Ԓ�?^O�A�F�Z-d�V�E��h���Ou�[$P+rŲ�v�655N� �H�P�YMA9º�ʸ9��q�����-���	T���_s����xa�n���z�ա�5�o�����ɡ�`���j��{UM����x��k�s�ߨ�i�@��?X�����`�d�!�I�ŖmN*oM�3gK,�
�E{:|@�a'��,�S�?!�*c�����$��!�������/�	�@���ޯH�����%��;i�g�d7�K}v�L�a���87�� ;}�*��l�����Cv��]M������ت�?T�����wC�\�J���f��KC�
���MY���t4F,����=Y�4���i��%��Q惧M�%!t���S~�����Xmv�Á�7���\B�E+�'���U%_�~��B�`�T#�(4��\��8Z�Wɳ�� ny�E��p]Ͱ49�@�p�E3ApҮ�-����%3����������4��[ϵ:�|��Z[<��)��(y��W
�S�T�W畝���&�n�9��z����m����p���v�������v:�Fʭ�������Y0"��$���T�_~U0�z"{Gwc;碚�t�ȗ�/��r��ث
��5���,m���ZWr�_��D����~>�-j�ؐ�Ө��	��'��PyՓ���<��xj��6�QB=���n�A��z0Հ]L��e?R�V�y�p�\�у��	{LKm�������V-�1�6��:�Ǻ��Hj��f��-���s�5��2�3�?���vk���s��g=l�5G3|���lW�B0G��P{�G��Ыm�_:a�ܦ�ߍ����)�K���g""�Y"BeR�Jٙ���}�!5ʖu"�(ْ#D�#;3#Yg�1����z������O�{����|�=�h@ɘ?�Q|��n��*��ĕ��w*ZNS`����::�Z�`&�fϘ䞌GK��@׹��%a��l�WY5�~XI�I��(��;��x(�T`�5�S�����Z�O�K�|R�^�É��q����
�-c����,i���QJ����O��B��_��5?^��T� ��w��?����5y�p���!���C�s�z�<��{ҧg���7X=o�/V�xs�����t��R�+"'[޹�XlL>�0� /�sn�y!�J��ٻ�4�}}���%�/^�a����|�_�;��+:u���������[����%�shlO���F���[��˖�d����3�̮G$�_��y u&"�⬃i�'\sE�����<Y�K/�
;X.�+7T�0bE��|�mؖ>w�1ӭ��m�o��Z��]�%�%S�	��{�^F�DbG���Ql�mN�k[��n��;�B�ofG��| ��T��c1I���W+����}���IfC 9�x��S��/9κ�oԪf�fd
˱��
X��Ň"�w����?�o+�?M��L�Yv�S� �؇
L�Ja���j<)��f����	��h,�����?(e`��Q���1\�,%��å������"KA�M�쥃���Zs垹�u�ep�	����Qi�ق��9&-��t�r�by�A�e�{��C�(Y���O�0��Z\K��,/,&��d~�d�k,���1ߔ��LY�J%�X7�7l}�"�[��(��G$4�ƒ{&=Gb��`����F��O�q=6zҝ&�^0K�P��|'�@�oIU��3�y��SW�Rz>��lJ���) W�O��0B�gaQ�'�L]gݱ���x�ѓ�n�W��������>�)���GqCE*t�?����Ε�Z��L��!{(짪}\c~�Ş8 ê��P�w�jw�p_��O��u�@��ӹƼ��|�\������뚍����$�p�|��Ɨ�� ����E���n��o1�th�7V!���,O^B{�9����*��E�*L+.�}�)NT�f����i���3e������D�Ϋð��&/{-I�d������2c��#AW/D�� �HzP=+�ve[[[��M��Y-���K���$�R�1���L
_�q�Y��`-8���Į��d���@�~Aǰӡ���x%,��]����T8IݺLθ(_������$���E�g�ޓ����+����(�h3������2�HXs����N��Njx�k߻z���E������:Xb d�.�gkM��3�v-VxƂ�g�4롬K��vx�͙�V$C���v�v���� r �c,/�ǟٮ���a�%k���{��ŗ�#��c.t�U��z�>9�� s:�a�j��E�ڶ>� #*pmuQ�w��r5�!Y�s���c�.�*����%�2�����Z�K�Jt����ޝ�N~���'ڭ���
b���!�9�o�PF�Ȗ�N��V�jS�bt'�˖��y���D~]̸��C��d�O�PxZd�N��sGft_���"����ڐc����R�EY�鵊o����ʻ�[Y��J/弅Iz��*��cw�c��CB�ֳ����3�֋`�ʅ��{{�I�Jƹs�<�9��n�|+�FG��y��v�����~W�e�u�n�p��*�<��i�M���#_�@?�[��)���_�2�@�AD�~%�q؂�3.!;��?L<��T��Me���i ��V:�����7��
Qj9]��\����w�:��s�X·7*��͔�������E³/),���8TI\���Y�	��@���,�p
�J����?<�E��?�I����	4�Q��ȯF�.U�rx�����/:���u���G�*b2��
��_��^��`_@��)��݆�y -.E�<%!K��dZ��?SlTZ�G+h-h�1z���E�1ʵ80/��<���V�BC��J$���GNCp�N�Eab���B�Ӆ���	��.���ýE�����pp�F8����5O\���󀕾4=2�B���J��3<�a�Ǯ�I���7��!d�h����X��olf/����"�<�bw�Et,���@��H���k\�L�x=C1ȩ0���p�>۸���lG��Fc`�K>��@Y�e��U�~{�l<�yyC�m���jw�D_���۫kR3��w��=#�CP�~�6d\���C/�7/�]>�`t��t���x��+I������Z?�7쒡�Q4n�`���R'~e��.�3m�EA��Mu�M�?�ľ�/�؅���Q|��A��/;���ݜebnC�V�4Ю�_OO�}�z��-.r��mW2��?�$}����-,��ǾeW����(��*=��>�BkͲ�ĵQQX���fO�=�檭��Kk� ����N��/~���親Rr�R7Ý[R6}Pܓ#|�k�lR�E;���~d��$�$n_�V�:v��YZLOawލ���G�T[��xTz�4O�g�#'�!ъ�-��?*e���Tl厯(������)|�f��u~eЖ�K�w�_�*a�D��1h�Xk@��cva�mZ�d�wK:�<��㯌]��/��+�wND��}ey���k���˿- b�ۭ:Q�+R�|�B���ƒ�W�]��9f}�n�U�"D��u�Y/�x��d�~�	P�gG���[�,K����̌g�$'���7���[���Շ!�z�0gM���#V�{���������Ô�MI�����nK^8hZ����r4�0����I�T��7�S�*s�=���^V��p/�P`G*<��m>1UF�Sz�>�pU1J���]�k�h�Б�pNm��Xj�`K���zα|`�W ��oa�\m���k��G����0��6�`�K�Y��uo3E#F�yJbb�=��%����UX� c���ʭ-_�|ݎ�l�k�����V/�K���4ٓ`�Wcy��M��&� Q�TU��\�}6 ����ڍ��$c���a������k���Q�o��m&�U7�}[�{��Jw�q�j	�4�9#u� �z?Y�<���nG�X��`�U�9��&�����E*��[�!��������nsB���ި��5���=�b��A�
��:�ur�f)�����X�S��'���H�� �-����VPK(d��`��Vi�{�ns&+��^��^�����镳���y1��>�o��W�~I�ŠȥG��C��	��wD�>O֞+�Ô��>�.jr�=��t6WjUڬ^�΂J��T��Y��^�^�]e���֨ADr4ˆ�G��� ���:zM��}EU\m+�WP\�ɯ4s���e]�\	� (�`+]+as�j���9���JP�<f�ԥ��;�:��+j�yn7.K_��c�D�ô��ع6'�����/�W��m4�/3�ڄ��	԰&��fZh��|�W ?���I�=�Λ�*��4L߫p�A0b�Ƥu[��͂�%@,`��3�����q�{�0Dߚ!=��QO4n�ݍ�>���m��D��$�C��v��g�Ä���p	1U��]�7��W+&�����B{�P����fI�� F"y�A�
��bW���;[ݨN	��$�>�v�� �%�˗D��E�z���	;h��* �y�Ɛ���.]��)��-/�ڶL�abh09�n���� �Ly�]�uԵ���|sR��P�ޔ�I"�����j.���V����?:	�q&p��A�4-}��L^���y��$���<��g0;���=��)���ޓ^�yP��ط-&켵��}�%睡��z�g>��i��Uz���;9��Nxi�[�����З�� ί4 ��b��6'��J������1��g�l0��.ǽ6�:�_��@���ez���.��57�}���Д��fHv��GeZ�ԏ���q�'�]0E��L˺��+��{q�"�f�I��K�|�4#vf��Hm�=��u�󨡖�r�p|�?�*��sºM3�O��&��U��#��R��L��������?x��)p�N�	[JW�b�L?<�l��C;;�r��������(�/s��+Ն7�]�u�]zz#�g�b����1?c>F:�i��`�l�ߕdv�e��4Q�>��F�f�ǌ�eF�C5�Wa�v� �TH\���͂��,蟝��\�i�CCڠ�E�u��{��
n��j�ih��s w�
��.���!3�1D?5�)�x�(����]������2�kAѪ�Lp�_]T���� �#���夒��ӞsR{�+L?����G�T�"aI���PQ; �zG ��8�/?�>����4;����S��4IAB��⮮�]��GՅ+~�]2�?������Z��,E�c����
���� ��Ժ$m��� X�pp�UV
�x�a>���
}��Ν��.9��ث��x�اAC�]�~��)~}����-���J���{����kH���A�'@ɫ=�(�D��A��ʝ��aR"xY�O���(y�E���}{�5ۃ�Q��Ĺ!���'�P6����@�+f�%V,dc��5	�:k2�4@�識��2s�>�����B�U�t!�|��F��K���C�G��&��N�_@R�f��GF�RO�G�|�\KNԺ�W}�W��B�9�s�7Ltuu���i?qB��є0�v7d'����x��{�P6�*�S�\h�����A��
�#;��V?`�����5&m������R��~E��'�o<� ]�w�3���2'�t23����n#���D��>��Ѱ�=B6���dt��gU�Q>צ�HBp��]�'K����ϏW0z�es��0uG Mߕ�	��HC:�ZU>����)���y?��\���d
�����/������E���L��卿<9��^�1�_��¾��T2/m�����q!
�|�e�nЙw���~�ўC�ұ,�X����c��sEBѧ�����we��W&�'�ٿ6�,���7{�����s:~��e���b�H�b���4�n\�,V�-����]�I-�}�m9Z�?T���D����qG�4�~&�?��-%S����>?L!ZD�$A�]�u��!1�����c[Ɯ�/��zg3YKsɜ���Tk/$y��
9po$~�)�]�t����x1�(���R�����s�ԄP�3݉�
�#�{(�)'$��2*Z�V�i1d�����5�sV&a�F����2��R��>���m�6I@����TL<.��(��$���uJ<pŐ(Tc(���D����+����t��{�4w3�y�[����c�LM�	�n���~��x�<�hr�Xޛ;�
�yp�	rz�Hv�7xy��l��f[!��p^
`я��}�����z�r�8XTT��\|lx�>�!:Ŏ�#��J�N*�F?�bP����Y�v�0�\�Z�]�2'3ܮ
:�\m;���f���6V�|MO:q:�
~:��*�a����#&��u���G�x�k�����EWѶ�R�]y����-N�!��v�p{A��!eMJ��N!᧶����-3����1�P\U\�}�7�'P�TT�j���h�rG���Ў���^��j,s��
>�7@=�w�>���2yk�\%�'��� �v��Q�fϪd��C�mf�1���>�����
�A�拢L���C�k�f&Nv�j"��;���g��7�,)MZ�:M��l��'��P�{ �ȇ�p!�r�������8�=�"�?�BΛu��\�8h�Y���\$�����G鯊	����Tz䲥���/"����V �����]'�nG��Oy��u�� �d�:��!�az�߶�6y5G��w%���f>4|ËmG?9�Q`G�A^�Av�ɼǉ\�=q�˜��'[Y���Iu��v�����]�/q?1���r+ �y����SV F� p�s�jDb��a��x�I��g d���%�격�{�_��]l��p�V���=\�_TM�M7un��)������*��7�ƹ�A�����%�h�/�D*I<���>�l�\�73^"gD�-s�ƸТ�A�!��0�[��QON��r@ve�$K�]��o���sQ��O]�p��+ ��N^�,��q���̜�O���
rOC��8����Ah�/]"Y�@�7��9����/�X �T�4�D��	��/1w���v5|�8� tiU}:9����T�H���$��6�c��:����2�����͎��Ds���e,J�W�f�E�J�u�K����a��w�ׯ��|��E>���֑|(��5��b�tT-JL�����^�gW�\�����U��d���t��V����ߴ�%�9պ��lڸ"���� �"�H�>hay@�dcƠ/]���qQ<n���us���ۭE3bB>g�\�� G�̕�{�x����y|��)� �=�'B'����k��1��R◡�������w,T�(�#"���gh����R�\jD�HʋXe�����������i�
���˪T��xpJKw ͵1�p�1���Q����fo5W��~0��x;�+��|~x�m�$�'US��Tp7�$��~�����X�����>8q����E��sИ6�!�>��ɧk
���`ߞ�%�����ޏ�#��
���8�q��vZJng}�9t&�Z��G�{\�9������#n}�;��J��Č	��癆n�%����Iy}w[|�N]b�tCm|ץU)�b}�x|O���G��ǟ��4�Z
i��0�=o�3}z�
�ΌV%��t�x_)�N�H!��[4�����?���W	�t�A�m�'�&��U��8=/q �d�����N���78�_:�����C����ͅ���ى�ma�Yg��T%OL�h�Z���d ��7R�M��$�����*Ҡ�����ڈ���E-1�xSXގp-��2���v�m�1� �S��a�(K
]`�-�}�E���*����QG$!N5v��vz�)�b>�q����18;���אe^�q]7ׯۥ�tv��h�U�$�=�E�8| ���!���_�ͮ�9�����-��w��$)H������.{j4�],E�'�"��;7�DP�M+5��gq��;r������A�mT���3��K`��q���F���
���V�i�?����l/��hT��M���Ă�L�R���L�("��J�5�%����-p[6�3^�l��ѣ,�r$v�����W��}����D�;4��]��[#E�nJN�&X�B��Fl�u��:�=��Ks����^��[�Z�m
�Yz��̯	`���W�j��{?�Pi�H���$ㅇh�6����8�..��n��^Ҭ�x�som8�����S�� 4�tcp�P�2�U������Ά������Tx�l]�"纝PQ�U�I�M|g���U|���}jhY졈�Q�R9vW��^'�W����H���S���B���S��(!�Ȕ��W2�]Q�� [͗,r6Qi�j����wg���
���R<��v(��[�Y�H4֘����5���1:5�d#|��:�+�O3�&���O��S�[����sHUrW���*6�i��ɹ������ʡ�k� ���&(6�q���GO�8��U�u=��X��~S���q�?��O���❴
;��m�ac����̿���a����41v.�P�48}@����\��F�=7�/E_r��1|sQ�a.�m��n[�k�K��g�z���|Z>![rq�>+���N�k�3b��B����-r*g�]�,<�܀�J��BX*��m(�?���OZjYvR����x�ΰ/ J�o|B�̧z������6�?�m��)f��r�\��w����L٬��Ƅ���%d۴>+��g��u/f$y��2���"�R�����C�Ї�O��v����^M��TGV�Z���k§���^(u{7s5��'�a�n����E�zG)F�O;�<uI|f4�� z7g�$�r�݉ʫ��7�=�;�۱�� �$�6��hss^�x9T�;��ᔄ��ѕ2�qC�Y��;}D�wǓJs������B���}H�)IY%)����K9�Jy�����A��a��@�l���i��JK�"�9�Qr�eyW���RR���呯��7����}jYk]XL�8��Vn�gCHyx���E��뵓��n�ā�e2U8W��d�2�����	d�M��j��iW�W~��֢CS 6$��gA��ЯʒE����3
5�7�l�-v��>CSXfX��f6/��,L~���e�ص���b�����3�[E�D�#�9ky]��i]���9����{i�lV��g9Q'��Wa/�`�W�6a���	�O��=%W�o���QӃ[2�J \�o6��[�N�_;C;�6xߎSν3����V����ñ����z���L�L[��"��ɢ6�����l'�����j �frn8���$
�^]4��Ua5��T,4�toO���1�ޒ�h%�����ר�Y�;k�xb�J��ͱ�/��lZ�--L�s2�{�WGD�Oέ������lT��`
��sܞ4��*����U����^�*���
�zZ��Aݖ�I�:);��X|#ݕe��}�c[�A�r����C���4�?���*�L�P(`RW�t��sA�?�%����VW����]P��ˊ�vWص�l�}-I?�J�n�Co����i�쨲�"�����O]�艏4Q�w�+M�󸐉<��}S��M*��ג�����[����vm�S��;jŁ6G�����h�>��WX�p�V;$4������T��6tUl����R:!L)�O�_��8v~T���T�I/.��3��N�w���((�^�85 t�6�L���=��@���|Z�?���=i�l�,Y��_[�?JIU�Æ�J�����tZz�-�V���1V�S���V��m	�~S�yj-wğv]�N^v��)�_��1��L������A=o�L3=��;&�)��U�H�A�~�e��P��&�̥��w��GØ�Gb	�����]Fr� �eK^�����v�U�mu��e�:�".\>/����E��^9�X�t�i� �(�=���v\(��#`���\(�����cY�n�T�uR;����yW·������:_�6JU�7��w-Q��eV�>W&��sǹF�R�zltu^�c�L?�۪LR�6����ø�V�Vmq�!緈f 4HC�V��Ш<w�*���:�zH�e�=ٖ�&�V�o�{��2do߈��<�6�+�*엩���հlь����x2��#�G���f��d� s�HR�w���R,��M5�u!���KՖ�M��},Et���l�'g7I�ѽ@l��b?}�/.��j��|q�0YurM�{��:�f�Ϲ����>�gw�*�9�0�02.1���n���F�X�@��	ӽ�4�x��EC�=�)a��~�n�?|�����\�-��`4���{��`=*��b���0�� -L?���۲
����C�Tp�@�����<SErc�]&,����R�k�Vz.��<�����*w�
�=��>���Vm��4����� hExt;�t������yH�Z�߇�d?mO�����a���G��\�0	�	�j+P-FjmC�F�8D�=1��m�������ESSΆ&�;>�Ҽ���\e��<��/z�kW���NT�F�U�(b��S����������	J/���)�Zk�sc
��������T��Ӧ�����@v�(N�����"Q�]-�}�h-v�y��	<O�%��o}
���@ݶ7�Kްy��l^�s�����K��=b��qM&�r7bE}56jD���$s�uD�ȧW��5�5d�]�\�[�ɸO�[�>BfG�<����{�dg����;��ww c{q�FF�Cʯ��cÞ���4x�o��r,�B�����XQ��]Q�lo���9�T'����.���'X}۬�$Ɖ�p��ĎJ�\P�7��:�z�$���gQg�E:�UT�(���|��X�w�E��o?��P�m8�E\|?D���9���?�p�v8��M� �k� ����/�N�),�"]�ȥ;6;fyś[r��I(�탌��s��g>�@�>���|�s�}��
��'e9T��� rP��j@(�	�ؠ�����& m�A����{����C�H��4^O�7�c���3����N:7�P�h ������D�DE�1@L�>\[b�|��d���m̀���mS���i9�@m�è ��-N\���e�@�����s��)h��Y7p���]�28��n]��M+P���|ξ�{�!�b���h��A'C�����[D�`=L=�15��|W�Y.�P�rO���d�bl�i�]�C7)ˌƫ���	P� � ��mJ���)Ѝ�`�ԩC���뻘��&}E��FV��c��R�m' c 4^F(��ʞA���R��Ԟm�p��Akd�#*Ǻ1�+P,y���������]���(d��)���E�d���d�� ʺ�rT����k\�J�g��`�̭�����<_:�S��筐`Ԡ��,�S5wR�X}����Wl��<��qS77�[���O��:��L�8 G_8>Z��Ym�jG�]�VpS%��,Gݦn��f�\��Y�݅|�	�զ(�OW��d)�ݰ�_�*+9S�n�,d��P��v�����LJ�K�ߩ�\�]e�;�= W!+���
-�玠���/^�������9�W��n����.zj�6��۞�M�ҎN(B�/-�w:N����R:��颎r@RI�l:�x�>�k��Q��|��}�E�����X�j�P7�mV)ˏ]l.3�7��|�yB&��F(B٣,E�9�m�;G��@�g��D;�٥����U�g�wؗ"�(=���(:@�6OO[U�0��U=��Ο��5W�ǒ�I�`�����,|��^�����P�&y \� Ŭ�v�츺s��Maz7�U�w݀S�P����� ��gT��P`	RcP��Ciex�Ɋ	q�y�x�pmn��|������A�A��34�J�S�"T+�Ys����b�ғ��e:�b[��M���P�j���~��Tg�W�8�ސ��k��p���ԴOk>/:L�	-v���#~j�����0ӏR�ڷ�j�R�T�\�6!�;����\��S��2@L��J*7���.��,����I2Ll��'�l��,Q.��d�v���c��8Ϧx�!��������j�K��F�5�e|�6�k���`
w8Զ�hU|�y9��ܯKN���@���^�F�R�W����ƱC�]�O@�)a����>
�*�*6u�V� ȾI@P�8.�
	-U���nVz	�,\�uK��RU�7��p���Ɗng��צ�hں�����'�Q:�o��	N�u5���s�s�����f��[��OW���;��.��
�{������ Z�Î���#�R59/�ގ*Ao�s�`u�S��Tx*�_:a� �oפ�ܰ5��*������e�j;/T��Uh;��x�c|�S�K����M�FBQi�oK�i%������?�~�m���]���-T�g~�?�d��Yv����)�aoG�_BR��f�*��͠�G��D�f���,�2��!%��yvopQ�sqP@�pͺ�)Fg���kf�H�s���P`Z�;�{�ߜ���:[&&(c��Z��:ږ"�P���'7���a�Ql��<����(���6��n���c ?e�����J��^v�S����M>����L��mJ� S��|�Ț�QW��mR��������r��]*��.�����3��,�ۛ�_.���O9�%s����eE��^̨����9:��r�Y/������-X�Bs�U�I���H��ky]ʍ�ù��q�0	g�c�U���,�������T�i+�S���nqM㘝�Z�����n�c��?�{�ͩ�w�PK   p�Xx[ǩ� ; /   images/628760d9-b837-48ba-be8e-acb7e191f55a.png\�XT]6������]
Jw7� ����CJ

��0"9��9�t�0����}����s]�5���Z�Z{��ޜXmMe�GT����T^)�FC���a��`���6�ՠ�ຽ2�DC3U��y@�*/��vw�� �痵��H����u^�5NhRD�k�9\�2��,{��s���Zx�C�'-�l�Q8��SRN�k9�+�V���-��_}=�����L�ρ�;o��<��=5;�Yл@N*��}�̚�>K����N��W�]���$1�:�3��B0�������Y_�l�����Y�GJ�a�Ǽ|> f�_(O���3@B �(U��r���~9 �IvkG;�#ZV�p���ę���'��;����5(8q}n�?r#������}>�=szTR��-m4y�L����߅H֩d.p��٫]A��vT���}�JFwu����O
��tbQ���2Q���bcx�y��'��"�l�'�"�,�Ѯ�5��Ճ3���Ͱ���y��H��C���bW8�j1ѷ�/�[���t
̏��������C4̔�g�]o^���������Geh�o]�]����Q���GY��ܮ+�
>N�aPv��c�����OL$���tDH�^{�ͨ��_�z�����Ge߷��7���c����[�lwIB�IK���
��oU����`f���=2��w��F�	h�i!8@T�pE�xN��*�4Ṉ�,L�&�����D�fi�oR]fũ����X�T��h�M��h�I���B`ɇ> ���6LT
����?�+0�<H��B��k������a��Q�C����DL��R/�>���OŴ?����u_"$N�������x���c69������L�c׬���$V�hk����} D�o�W����̛����mA��	o�eVd�k:Y�sM��;����OΚ�c� 6��C��� �h�Hb#����8z�$��uӛ)��m�11AxG�T��ޠ���-{�GtK#�m��x�� �^V��TU��F0�7�z�ˬ S��S�"������?��n�~��0<b!Ϛ�Wi E�.1�SG�g�$	z�q�JnM�n&�J��@\/ҟ��#������hO���I���_��yo/uqG2�A��Wg�s������h�$5�t���\e~Dm�c2ǖ���	�ta�S�[��>����"����[�v�IῈ&$�v�tӣ�������N��9��æ�q��b�H>�ٚ��߬��-�Č�VP�tm$�s�^�Z�ܺi&e{ї�h6�����]`
�o�F�<\��A0�RL���/�\a�? �y]-�-4��G�Ujg���{ah�ϱFv{�O[o��c�[=ߕ*)�ٍ�>@��7P��r�e
��2(�8`��Q��EFQ��i�ꕏ�_/f����a\flʯW�&q�j�DJ��Y/��/غ�G^���s!P��#�Z+ފ�SW-���'�O���*�M���ڀ��<���`���H�hd�iy�/���J_FGxgO�d:�!�q�z!r�4s��i*�>�R	��Mױ��q7�fKs}��[�9sF������Oē���F�vG��P�B(��Ѱ/d�!�)�H랯��P}�����,,f@�k���CN��s��B���Q��x�.���B�@jM-�3D����6:b,^Wk	�[z�@6c���v��2�ڟ���C���+�V>��N�qr�x��&�σ.���F	���C���'g';qp��6�~��{w��iT����O��X���դ��3aࣤKj�p�8GZs[ �P<~�9W�?S�'������i���궛x���|-���qg+d�lz6(T]~:]����������7^-����|� 72 9B�0�� B�W`֌(�Dȗ�M����_��ړ>߽%wRiY4^�T/X@ޚ�$�}��Zm�J5%9_��yۓ�d�#O�����ӖaO)�~3�Ԃ����C kހ-8�P�9���i��0]YS�Ez;�[g0�7׶Ĵ������𔯀���ȁ�8Bz�w�@F �~���������GVqd��!j���)�sJ���K�w��oG$0���k̤ �<�?n��1x��3�}�8a�ί�%N	#i�������-�h=�Y^�+��|�2�XC/UdI��3��r��⣥W�����b�ȶ�������I��_��J۫����RBв�%�vr��R|`LzV�jy�;�\�e�)��g���d��o���]�MI�Ť�{����R-�؈�]�w�7_C�����G�<�ޙK`:zR��!�.�l�~�����&��ELqKD��rTT�d_&���������Y�������>�k:F��K��B��Kddd�����쪀K#u�Õ�v�Tfv�C�,^).�n�C��G[��ۓVZ�#��J*�gX�Q���-V��hk�]�H- �F�rraZ���������#I��U��D����!�x�w�I{/^�����^��}���r}s��[��q6��9�"Ѓ6)%�ʔ��#�a��j��j���N���V�ӳ��,gu7� osw]h>9&��~�{p�-p[)�xi�Y�|�gY�]������}�=�k�7���qk�w���_"yyk+:�T�bJ{�UFQXX�̖�56��5�Y`s�0:;7O���7�XX�(Rc.����S�9h)F���I�#(��$H�-�266v#I����+� Tʋ_�WXR׌�����;�� `֊��i>>Շ�,�!�!��� � sPD�����V5�h.j\�7� Q.���WaY7�>+���<����Yixh�ް���_mG��}(+�[��s��RM�\������1�mY��}�#�W	�u�~_�զ2���
�(�����е~>ِBEQ�/!*����.����t����:7gԏ���UU��J�%hX3{��br�0˘�fY�ۣ%�����+{��D��>aIؗ�l��y����>�h,'p��5�f��R�r�0z�MoE���~j��hnz~��H-#?x�2qWE[��+�↰l�ɋXxZ�7oa�la+�{�f���4�.
�/�=ht����"��u~��T'=/ѽ��_HK���Ғ(;)$�F��v����;y��ŷ�^�	
I�c����s�4'p��� Άz9��� 1�<4���Fxj�3�&�G<q��3DZt6@v�s��t�Q���C�̡3qP�A$�(E=Y�r?1�6�JAg���Vb q��Mɓ�x�w�������z��h�.ɦӛv�̴�36j��kJ�6.��F��4w]���l䞭�Q߂f��<�JK
���^9Ob��^��%cW
K]io.�~���5oh\�*h���a#Q%E��#8!���j�y���Y!~��_3[��ڗ��,�9����Z��m�ͽ�{2$����p}���h�����eX�l�h��Fk��+ÈR�C_�M;&P|���(u��a\�h׀�js,���U-Vk�ʑ��!+�nNW�D�ҷ*C����Lf�
Q�dF�g�˯k�Bx�n��PA���K`�z4}��y�h��4P� ����rC��ދ"m͉-���Xlp$?��:����n�p-G^Cnv����������l��kC�6#[+*VU��(�Ѭ�Q>���Z��hu � t�0�Z����l��zՏ��}2���;UЉ���H��"�	6�0���/�����}���2��� ¼�m{��p��,�]�����[΢�]�����T�3�:о H�O��s�>��k�Ís���J��n�Vw�n���z����7�厲�������R�My� �;Za��'������ko�
�1�;~Ⱦ�3�y�vK�L�Z����u�����-����*�FN^cژK�&cILd�bm��7��2
��;sF-4d�P4,���	���d<�^8PRW)�(��:��qI[ ���Mp���9G_���4�РPI�7�_�2�����Qlo���5�D ��'�#���D�[1{�2_��Gs�OUR�-��Z`��zR��H}�Ō#a%:�\�%#�@�ݑ)��w������acT2|�]��˲1�2��5TaY���P�x(�V��WTĲH=T��E�oD���*^��]?���F�+�ϝq��t-�Kv��uůs.���D����X�H��~#��~+&�`��ɳ&)I��'��,�`M�jE5k��I|t��eH��؏��x�����k���\��6�_��~(L�-��ĊW��N�����q ���\�z�@jfh�D�?�͈lgG��g��g�y�;�O2l��Wd��#�$������,�^�4�� ��9;u`���p�4���CU��Ǵ(.M���^c%��,��b�b�b�6S����Bs�y��4x��"go�����
�����ȣd�0���/]2������k����ż� l/���6���>5��,��}�Ua���\�V��q]C���Ϝȋ%j���o�+� jAL�dY�%H;�̳�Dwɽ�H��gF*���{s
�'�!��@ �g���0�x��p�\(�����=���2�?�t�a�:[��������q�(H:���hN��r8 ~�q�m �k���"�`a�%`OF��O��x'��i��R�]nrOɨ��2��'覯[�X	�K�Ru'�Y},o����9(A�V���K�b{��S�4�Y&mM�36>Z@gr�yy^��k��ׇ��\��|�cUTLG^m�m�*4����Ӧ��d����rk�V���^ꆌ����5!�����P��^z.�x�ܿ0R$J�:���L���o��X=M���]�2��k:��"u>�zZ�cl�~�e��"�A������	��+��ɝ�M��<�$2�_�E�-d���I��ţ�za&�_�����z##ˉ�������2������Yc�âWQ	:���L�%�Gs��&o�����į^M��mZ����s����$�gA��N�W��DC> .~���a'Kۍ�r(N~��'��ת�{����8G옳(+1��}��&h��$�++��`���J�����jD��N�O˸e;���ʎ�ϭ?��P9L���8�8��'�ݏ1�ar����c����"�)����<Չ[���?��R^��f�z�����@��v�;ͳ=Y��D���_vvNi%��o�������o�ݞ�3����]}��JF��|�0���Z�t�>@ޖ��������[� ˿z��&Jz�_��?��T���2r��`�����*�/P���[�2哌^͕�qK�F���߃��ٓ+�7?\=�0�����սY��I������<�?� �.i�z�3�R?��N��M� ��Dڏ�-e-��|ɍ��r����3U�Y�y�0�2�6sI,=Vw���3U�������y���Wix�4
���{��
5�+�p!(X+��r�M~7�O����m�<�'��b�31��f�
H�4[��ǈ�`����2Y�ٻDI.�} ����+�@�F{Q�W��]]�W�.������sW�ոO-!w��_0��k���	������X�D\2G�S���Ovh2��j�=�L����.��&��m��]�=��N�������!2룥��7��H���܄���bf�/c*T'a�y���0���W�j���]��DL��I'�|���j��(1%9vAŸ`��e��Q{���i�;>p����@x��
1q��a�f[���ј
9��G+�;ޔ�P��Z�Ĕ8��I��k�߯��b�W5�PL�3b
��BoZm_�~|e���e���3�q���NH��ŗ�)(+�?���'囩Q,���\� %�:����짷�����7.P
K��l����_;N�x�WD�®�\���!������f���͒�_5n>��Ū���X���h�;BW�$���S��Q�����+�ʍ4I@R"N^�\j�ߔ��=�!�cNS?}������(w��ٞs���x�hT{#�~��@���Fږ�%���wMǰ�PQW?�o˞#�7U�RO�Ѥ�[(�����ќ�G���b6Ue<�=vгf������x�y��x1�pǜ�6C�6���n��B���!4��,)7;�����v�DR�x}��6���5%���t^?Y@b0�;�Mq!�/9%�4��T��
ivt�����sPk���g@���n��j����~� C��黺��0_�z���.a(��q�y���U���ܼ%@�P��2�nr?�v^��*Rxd����c,��T�
Ӯ��J�]'��l��R�SxŨ_g�`��O1��j/p���\A�[PYY��,�����zsL�㡤�k�>p�����8�er���#|3˳�����z�xunE�3\�MDd���D���'��i��o}0�8x��-C����)⵭�y�l�6���r����18���}0N�n��G�\��c$J��7o��jWR��W��c2�%�8ݒ��� ���L1�L��0r�y�1�\�UX>�T�R���f�G"��$x�����7yP�;�*�+����]�sT�P�k�'Jc��Q����`�q���^�ܙ���	|�m,QW�0����.y�iѾ����?$��?"��R��-�৬p^V������Ѓ2;ła�⨼aD�CM}w7q��R^��{�uD��[_��M�0�1~AŤ�&�N��C�;����*��S��úWA?�����@���ӝ!�5HGC�D����n'Q��8c�g�Z�A{��55�7������ϐ�,aN�H��G0ڠt"?Q-o��ޜ(�A��č<bg=T�)�P���[Іj�G>ȡ|�q��rk��A����~�B߽���d�F���g�N0�zx��^�(�7Ӣ�J��#�}6�q�d�B�z��/J 2����8J�88-�<J:Q�͓"�����qx�c"L�>(��/�c�F�X�$!)F^G�q4��lKZ� ,��y"(/�$L J�T��z��	ep89�2ޏ�Q���/�`(2�ZTߺ��ΏR\�oS�"9���a=��죶���U�2ʃ
��C�?�h־�V�6�FQ�l�3�Q�f�XK�b��Z�G��~���{XѬm��,�Ȍ(n������ײ\������\�{�Я�r�[��*�{~�6�=��Js�)z����>��`�v�����k'�ͤ(�<��QV��C6�~�إ�l@l�*C����7���Σ�g� ��h�ྱ�K�����ᙤ�'X淏B�Ƶ]8Z�� �o�7�!�>�?�v�p}�9���Iŭ^&���7����3��R�Ԍ���kE�N��>&�V�dz�ޝ��RIf���-6���9
ш�^�~%�l�B<V���u��4n+f�Q	����tݦYc�u)��˚���	�}x3h��5(+7�?��L����=��~�-���=��|l~��Pӕ	
���~˙��ٴ��TTPJ���!
�C�Y�uPJQ
%Z�*�&q���)�U US�9�qaI�zX�+�j{o��T[\ǈBԯI�&Ew�����Q�������b?��b�_w� �ڳ�KK[8k�'"9%ϑ�j��@3�������]�h�n� |���<��/�B����((H,�^�5���H�n�R�O, �Y� �
wi��W�:�|-��7��=��`�P���?��9_ճ7�a�����*~�rq� ���1���y[��2�ei�Z}����k��� �M�L(*Iz�t��8�a@��1C��~Om�@�@�l$�5�ļ���izTk^0�*P��P��ع6��Z;�SS��ݎ�ѥ$�o��o���o��{ՠ��cΡay۠3\ϋ��%S����m?{1:���FQR6u��9v����_�RA�*�߻�v�\�a�"I������+'M[6�u�GP۟9<����7_��h<Ql��{���9��W�����Ϩo����%Xw2���!.�?olL��ئY%%�&�)f��2�'oN�_�b�^������0�~��*Áu⵿�o^�a��:X��/+zv�b���p1���v.�Kt�mYN��^21��q�� ;*M��^�ӕ+U���L8^۳/��5�kLj��3����]?޶��o�۝cK

d�ߘ�����`����h+[�jj�������/�]LL�]���m"<��Y(mUҲ���2ǰM�!}P��r�����~������W(Ev��6�󶌂z\�f��w2P����9�E��Kk�����$�<�ˎ۞J����rM���Ȭ��������U<@o�[h�x��6�s��i�f�ώ�싙���"͵��Q��e;_p|<��D�h��x��V��E����kO��so\����d�X!����s?��
�[��a���F��Z+-�}k��H��d�SM���ڏw���� �
�����#eJ`�L����$zpI�ňc����ѻ��l磓�|Egպ� ^������ZEZ����&M��F~�]PQ��n�B3�^E^�,n����~�<xDu���z�i���	%��O�fR��x�����Gܞ�P@�M%�0A��JP7��}�/S���T�FP:j�G`1��Y���H��)Z�_o��7������ۃ�I�����;>Hj����3Q��R��@��֦z�q�& �uH/�f��W�dᅕ'XMx_?�Ʃ�wp%`�=e�YSp�n�ˆ�t�L��Wc�������6�Kӭ��3��i��Uo���_�M�Ь�gd��ڂ�Qn��Q�"�r���T�~&j�Ws?q�X�PUm�,/g�;�.iq�Tk�M��7e��:��ͪO֘�kD��M���D�=��77�(�a� �V���9sD]ad���n� _�ZNt����T�+��}b�%��@1 
��;���k{�����v���g�(�)eܐ%�Mߥ6�<j`w����Z�b�&pw�t�uS���r�n��@*�S��؂�BE���5m��
��7�;��c�{����%ArB��������.tYߠvƀ#]ڛ������E*��3_�����X����g�&��_�I���pR���y����Q%"o�RTPǏ�/�ut
����+��=�#���z>��xAD��eo.6��������8^7c+]�!r���g[fF�;����M��xL��^�\&a��Tiv�~������خl�P]�t>��P�l�5�kŇ��f{�K&���)�k $jxùl��>�:��^k�0�kJ�0�����ʼ@q�����ҊD֖��]��'�kG~�b�4*H��ƺ���
��Eu~�+�D����a���H���}_Ț>J�3OЅl�2�?=U΋�P�{}�t��O�ߥ���;n���k��L�@I�׻3��T=6��O}歜Z�k��Z��*~*�j�5�9�阖-.S]Hjg�%M�G6}��\�S�����iU}^�)��=�\[��]�=]-���f����8�};���n��ߗy�{P �G�Xn���)��ǩ�(ՠ���T-�߯��^[K!p�g�ESPT�;�r��(6�����5������b�RO�I�ٲ���T��K�艊���u�rZ���J�K JwA�!�0��|��x��uF���xwC���n��*^��f���6��P��M��y����uܕ"���cm��<�}��U������K�j;K�s5�~����۶Ń>d#4a9 nyz�����D�O
��x�$9���Dl//�^֘JC���	Tt�jZ�r=v�2]z�����WJ
���crWZ�Ŀ���H#cJ�Vn���W"��;����(,5����O�"D�?s�3޽�Az��e��L^��5ɨAj, ��~�����Ze�]�=!��᣶�k��)�<*i�DJ�n޳�������M�1RMU��]Bf@�9� Y}aT�E6օvO",J)�"�(�ߘ+��'g�F�L-T��u����ҽ2����l��5ׄ�!���G��ϵ9s��s���J��%����<p� ��'���n���˶�#��<�>�-��F�\�s�iH�d�Z2R�!zJO^J�����A%��)CX�0��ַ}���v�u2��wY7�ٚ�t��3������fO.�mq�"Ra�M�(Of��<�>�Į_�H�[j��I�=g(vY� j�:��o �xm;������]��G�M2TȺ�Y@�1�!�"##wo��g��5�}X�Q��p1]��q٩I����9C�	rJ/P���[�a}Ӝ�)���@\�e�����T�piI"��;�T-��=�}��%�nu-޻%J0?�>.룱��-KǞ��پ��*|N5s�J��
-�$<�kD�C_�Uw�����U���"�6s��N}Gg�L��A'�ƕ)[��%������t�oie�5|ك@տ�jPeYjΐ~?v�t(�Ӓ*��G��/��{<����t r���0���;
>a��6##"֙V�P��S3{�QY�����q�״�r?�y��7#4׌Z��JA�������& *�iY�LL@��S	����*qbψ�f�MY�\ӗ;{�Q ߩ���Z���ӨEP+���WlEq�bH��\q5� q7�R,ۻ�:%�dHw���\?�KNYz��pā+��KM�e,y q+�P��Sԭ�����r����MLI����%��
��II�9�>Z��]��؂E&oNu�[Js�O�F#����a�º=[I�C}��)��NÕ6�l����'�l�F2�x����W]��yK?��4k�	
���{����/�Sȕ�{`{��U�E,�Q���fAȽR`-Ѥ��9�5�;�fQ�
?��yB�o�{%ze}��`|ڹ�T���K�T�����}��G�oTA���Rܦ
El�d@�'R&��G�8H�U=��6ʓ�E���]|����'0�b��1Iɀ�2 ַ6v��p���x�tSip\�����-��U8����(�ܨ4�s�+��=��?{BA�K#�J���Bׯ����N~NOI|���#A�P7���Vg�.� շ��?����c�H�2翙L�F����v��}4���B}L�˪ݖ7�f���n�����74�Ag�Y�aCR��7�_�*�9�% kx.y���Z��~�FL&3?��Z'ԧ@����M�ydx#�yƃ��ax�ﯽ�Wj1x�9��>�5O��QZ�sDUq�ɢŵ]�.��;����S��Js3�� "���fDe�j�\�;��*���vҢ$�^3��_1�@����a�eot*W�����]�:�$�\�oR:ᙊ9�M$I���	���d�l���s#M�^V�U����nr;e%�.m���?��ԕ3���@M(>�7w��CQ;p�@�������Ak���k���h�˄V�A��h�2+���e�j"FP��.ۻ�˓b���@X�D�L�Jɪ�̵ֹ�1��&qY�W�y�Jخ��gn𥎩��ȃy�͖�mGۯ��ZȆ���QY	�Z�7z�lk��9m�uP�l���!.�-H8��g8�&к�'����El�ʆG󴘾G���HqZ���ȝԷ/��v&�1!	;� 0��fMh���n����ύ>{ND3�w\�Sk��87<�zBn��E�4�2���\J��՟�7��_��>��&d�h��[;w����V���'T��j>�����E{�խT�zH9���k�|HEo�kf����aѢ�v����5�l��~���1��>T7��>�:���Sߟw�L�#���V{�8����ڏL3pN"Mgco�eJR����&�����#������;�Ԕ_a��'sl�3z�
i�@�Z�y<4l�݉ҥ	�x֩�J������G�;�
�@ZR�fJL��d�F���RK�r�`������P}1�N�:|�D{���"u�{��:�(%�~�!	�;⯵����[�H��N��5i��'��ڟ���N��9��Ei�G�\ۢ����	�Fi�O_֞km�I�kZ���\���m=��+ʵ�Z<��YE�{�g��
���JW!�u�V��������&-�$М�1-�?�~�͑�z51&�<_`^Y�>9��3$�k��O�G^�)��Bh�*�Bu���(j�=$\�������6h)r��/��&"�j�z�����өTb>[��t������6*���<��^BL)�r6�v*��粿��?X(4l�w7(�ϺU\p������^�bd��P�~��Bw��PZ�j��ߧQ��<���*d�3\Iy^�����
:gDXo]����d)Qm��Ax�.�_��ѷ%�cK�]7�J!��d�!yh�	4�����Zw��>;P٘Z�$�1��3�f(��E�����;����R�ex���$�L4])�1�J�����޵5�ԨU�T�ׁ��X��W�jn�CE���~s�{���.�n)/�����L�$���������Qi�Wǌ7fa�2��>�v���1���Z�|NGY�h�F�D��#�nP�&�4���D4�u���t�<��H�Es�K�)G\6_l�L,:Q7��W����Ӎ�wm*,Q��z6�䢼}#V��5��Ĵ* 1UBk�@k��ۅ"C��&���DW&�^��h�q;�s۵��LJխ/��,��[��Ek�ߢȄW�T����}�������t��r�T���%s���4���qL�T*-o �PCsZ�v����jI�e����qr���0l_�`\�Ko�f�����[$��	5�_���CH�;��FW���%��?-xO��;-��O*V��ii?/����	gֈ�Ǹڿ:S�έ˯N��2]p�X�Ѵ����\#y���T����ٯ�I��9�
7���ך����)��;7�a�Or�m��-�nʶڎ����vz�8NOf-��f���O(c߀�� *ܟ�'iem�Qd'�V58�?Dָ[[�%_ �u����1��5�&z	"c�s��$�ӄ&�S=`j���bC��[ʭć�FPt�!�ña��2�J��l��LėN~OJe�I$��%7S���"�g�	Y ��O�
�t�^�*l�ȗ7J��gWY1J��R�r��Qu�,^K��]M�q'|A� ��T�0�8/��Z���mr��<TK�=6]�В��f��(���:�C�sߞ��'_��������1h��L|R��X�]�۫�ݻ�G�n��|���$��s6ix�w�v��-H��ڠ[�ǐ
�����nv�g�DI+�]�� �$�5�����Lг�-Zm:*���gs��צJaAwgv��Յp�3������3G'�<�'�I����K��1O(\��uD�c�D�3c�M���A�	��&�vp��f	Шr�5?�Y,,�6��~�\<N����ǅN�dm=`��{��?r���8]�e>n?K~�>Y�w�8��l�H�r�ɝ�@=	������WMU@���^��/�����릶篆7-4%��oc>�K��v��+�����Y?bt<8��m}F��3�U�@Ѱ�����m�����m1�Ю؞���oG��{�ߪ��9%% ~��ٖ��Ȍ�5Q)Ή�Uz�)�����sw%��f�l�c_W�Uf[a��nk��kל5���M�\������c>���-9L�7~H�mC K��MJ�=�J�]��R��xh�3Ol\�+y�y?I�e���Sv��@�Q��1��&ǟ *���/�u�~^�R"����n�6�Cr�8Ow�
���c|�d��*U�.�g�WŤ&p�=G��+��WgzG|��?���4�JB��o*a4uIM���g��K�i��*�����0Hr���ŁC�sV�4�I�#�a6��5�yq�U�x��ug����f�'b�b�y�E�Q�L��=3Ri������I�!���ҁf�\�󤱱���R�W��cއ�;�=l�3�3�s!����G���)O\��1�1��J	¸F٪b��ۓ��t��ؗ��B����ޏSͲ	��M�c�[�汔,=ra���(�PRT���{oJ'[�HGR���+��w�yq"����b��@yz�^d����j%�\���1m��B)��������)��_�!7O!�^||���c���	R�U��]��k���ոi~�U�J��ryr ���2A�,��!V��:� 	��m��jZiTWk���;s�E����Zb�ڨ���:�����1��l�6z����G;Lr��Ti/��Y#��7Wb��p��G�T��L�K����-���:Vр�2k+^��V��sv���g	{�/��WC҄W�m�~o�v�H�D~!?�]2�d�	��EP�-��ѡ\"�[6���'`�aҪ��C֭�����^�/���K���ƓN��B�}i����Zz5=�#����]_�F�,�	��v-�f���%�^��޲`�pUe��Z���U�֚ͬ��H���,�ɔ��6`f��WRC8�����@� t��Qs!椦�a4Ѩ�=zo��0����1(�H9�ƶ"9��,@R�a/J�n?R���fky�����
l��ޢ�ş� �nw�r�VU�D�R=cn����3ӢA���KVm�(�^�p6+�G���p�L��։�m�T?����Z������'��_�G����uLLY 7�4��D��C���!�<v��4�����G'��H�lw�_�R�D~�	?
j�k���PY۬/ z?~��d��S��R�J��F�y� ^�����lM�Ԩ0��l��H�N�+x��,^YA_���/�Z�HS�0=���QU��i�c�jI�	�g���{����y((�g0�m��Æ'�Gꪬ]~��^[�K�Q�m����5;�$k�ؠ�{��lo^M��9H��QVu�qoxP��/>��tP,+K�:��i#ٳ���4�P)0x`vto�|����+���!��u�ˣ��ΐ��ߡ���7ȩ��������k��'1j���[�i�7맟9���3��5����kh�W��^����7����G|��_/H�Sn�4�	�@�(ŧo%MZ�W�rŢ��� �<�h��L�1Y//M�u�,-�]���v��~�	J���<6�� ��F��)��L�

(}�sزæ�#EkŮ����0��uj���OJ2���h�pC��~M�[c��mY�<,?�TC�H[���}�=����QHlW��k{��&\o����ʛ�:5R�L�Ϡ�V������J�wsk�S�u7��"�p)=f���ֲ7)���D��o�`*agM�Ɍ��Ѯ58����Wk�g�ُ8I���-�4e]��MH�7�����vI�c�b�J�ʴ�W0C����[���,W���ZH6�F�H��
\�����hz�<��`Z:�S�k�'Ё�(L�:{���Y��s���;#��T�;��a�.�^i�g�]�ڑp�j�n�8ߙx�n3�̴ey)��A������]c�~���
�����7�$|#J?�����b0�7)���nQ���YƝ�~�}�7�i<"�k��mJ_h�%�<���j��|5��=/�s&~�[82��Eu���H���ȼ�$�:_��P��_�KZ�����Y���Qi,b��p�۸���qٞ��*5T�]k��8N�V��a�I���*I��.���[���N�_g��x`6eJ�]������v�A��A{w�Sj5�W2�R�T��Ĺ�Ĳ�B�.�\����Ԉ�r���4����l���>�?~�FE[���]�
�7%$�fIk�I{����|O��Rζ~����G�)��R�^��+����d�p��%���WG3կg�&NVD��9��{�J0yEI[��(��F��׸w¦�t�}���B�J:vK�L�=�`;�c��*�i��]�������Җfb�Ex�n�̩K�Y��3��c�ғ�"u�$G�(Xv��_Z(Dџ!�''ӵ�y�����C:Q�c�ܲ���r[�P=k������>E�����`�Э!AG=?��`��E��\�pբҫ�1�b(�j
��㛞V�Tw��-�rZ�T�v��@.�Y��ތ唖t����~|�uN�?��H���)��K����M���jL�ˉ��V%[k%��J�9gUI2=��KW��oӍ�4��c�,���g2&>�w�.�Bu7���`�^�:�Th*.�u�Ax���@�.ŋ�w��$U��U���R�g�8Ք�ۏ7�(no[�lLg�S"L+�8�&��O~a_ZN�3���*d$�D�$��"Պ���a�?���������5a�%J��ڶ��p��sm~�n8$!��k��t�!���\Q���������|�6�:���_~+�?

8�kP�B9�2��S�wշ�A[�<�5HA�v�;��-t76�E��M�ifM�	-�\�����%Xڦ�ա�}��ڃ7G��l�������|~95xA�iF=��n�ؔ�"��I�Ց��� �o��ˬ�G]�m˫���-~u��c�9V�AΉ�b򈕱�i%�Ѿ���O���Џ�`����#��fR�w.�5�����%ք^̚�o��b�xgi?$ԼcC<�<���}�q(	<E���L�����z��Ͼ�yc��\��YL͔��/��������H������_~=E��og�x���_^"O����?��2,�h�V�P��I�f ������;�f�n�P`h��cf���9�y?��.��ޱ~����F�bH�����Y��	�|lWt��U�;X�պw�*���]u:Ϟ�f�>����K	16���	/�B���]���r��«N��)��L&9[��^h����Cy���|�79���DF׽W�"O�L��k����:S#/ea���y$�z[� �0<o*�VV���#O�j�Ï�S�j�dШ�X6��(�qcR��#�P������m�I4ce�j;+(`�^Q�vo�d���DK�b��Ǜg`�����,�غ��R'��z��Z���z��6����i��g����L�ky��ۍ�lbD�n�5�48u¡��޿��y�}ޢW�1;%�gG��Nt?��Eܭa]��k�MqZ%�o�Tj7�A��&d�/��X-4��8�JbҺ��E���,8�NcUܞwg@���4A��;0���-bl�є�n_���G��?C� ��TSQ�h
�}Snj��5���5�M����Y�U"wJ��_x�)\y�֌��$�A�=��F��{y����!đ��L���?�j���R*1��:|qJ�~&E�J>�t����`
Ʀwz��Z���I��(�_�+��^���i�HF6�y&>�Op�z�?�OBL[,��쫟ڥ類D��zr��|,�cQ%$ 5ֳj�!��E=���d����/�̭f�6��4e�ɜk����~���U����dB^�r��~䴹�R�q����D�i��H�#I�g�͝y�����Ѣ�����6�t���� ���,ѩ9��?�e�0�x�\�h������ ���ω��r�^x
q\G=�	�{���ͤ�Ö�K�a�r����d:7���FĳTK{Vpd4�,�U�b��������V9�S4�ԧ�*F�SSN�D/�ث��H����F�-����5����v�L�t�Ұ>+yX*��D���{�xB�xT�d��ێ7|��ܽ��oZO{�z��=!#+��0�8�t�Kb�n�����V	��k4��`����+��&h�pq!WzY^y�	�^��*�M�d�dؚyt��&��[���ٱ�^jd:.D[��WȧR�]خ�/�,Dc6w�[��;�|�iu�)+�Խ � g���Ũ�Ĩ�أ�	�U㋧�vz�K��T�yE^B���q��/��	5c*��Фx���9��X��&_�x������W�A���6��%�q_ɱ|׸��\쮬��14_���b�9�}k��A���#�Xr�b� Ѡ�y���Cc�WiY������{긹e/�IQ��79ig��<�`{k~�c�4>���ӷ�����ZGr֋yȬ\F\���<��d����N$�םR또�9U�R�VaO^�J� B�#��9�WTU�EE�*D���<��~ac=U_j��09H��(�}�gt����u�������h:P��m.��|�O:���#>�$^����S����nea��_��]	>��7A���޲;�ݝ��a���ᩕ��`�)x�h�4�U���=���e���A�=<��Za1�%h���#d�t��s�������Qc�� ���M�X݃؇���`!3�H�V$��:��i�L֪�Xh�Y7 �E�\�@3z��uT�8��-,�M�������X�p�t����<m�89!�:V[˫�[Ç�%���j�{Q�ɟq�������^�|�Hgؑ>�$�B�ŷ�W�4zV������j���)Y�k��z�9WZ
	.d�gs��������4X�sp�m��?	n0[�S+�à������ꗃn�*�t[���� j ��HͲɈ4@�e)��-����5y��d=�<�H���;��~�=+5�
����-x�ܺ���>�h`R�f����i�X{�\���qq�sI�`�O]&N/IuN6�')�O0"���ҧx�$_E�˦|`�;�>^o���)��f��?"�T�s�8�5�9�EA$���*G�0v��T�S�
��<p������$HOݫ�N�E�ėV����ui��� k�����ٰ�ɧ��?���$�`I��>}/x����}�S~��s��M�
ǥȄ�}{3��$�D��1x5|��|Uo���
hނƂ�4J���6�}��٥�Ҳ�̚nb#�Ze�Ky���9]��/�7#F9߉��Bl�3��5u��}oRl�^iZ�K�c�1��d8�	����n{]�	q7����)���Pb�o��� `u��4!A�E0Q���}ϯ<�lqV��_<�s������.�[�I�M���N0�u����	�%#""6!�q���[�n�Ӛ�)��`Q��	���l��nYt\�;���d{���₏�Oѹg�`����{w|�zd��.KI��(�pF��դD��B�]��1���@T��Dg|vv�d�5�BY@V��Wo���,,��TЉ�p@/	,�&P�>��h5_���H�j����W�g���v�_�+9�gV��4�n%�M&�����x�B�5��.nJc��c�Uzh�������`����z��W��x!
 N_�Pâ��A���]��Az�1�:cD?@�� ���A�v�2�.���o�v�*����n�I�H���ջ�Z���.��6;�n�y1�<U�zY;�|P�Z�o��^�^F�{�̡[�$��dLr1q�,Q>ͫS�*���.�Yo?��E!,<&$��4t."�����U�V֏S߉X8���:7��i�{V��������T�J��B"D���i�Drc�b��/&��~�S�������(O�S��@���C�s�6��]���k���I��.L_��"d˂�(K�m�_��_��d�64	�~*j:��U�;��Z|���8�A��s�	x�'��G��g~��T���A/�M���eض>|ŉ$~��1��W;�"�΢"W��Eٰ`8ty��
�tV^�F0�`i']�F��j^��zrp�c+Z���A�d������Ӫ��v�34��D��7�}��U�VG�Z�%DV�g#��Ks�����vn���&��,�� P�߆$S�����1��ͤB�I��C��2�j��9�zê���d�Xp�^��l)/t�îͮ+Q7��+<��Ѥ=^ǟ���KC��Ym8�vy�g��?-��m�{��ܶU����!�Ȯ�^+�Oe*4 #{�SBn�u�7����f�&-i����SeKx*��O�w��:̲=]7Me�o`xO&r{*�]�����3��c�g�S^"h���g�*��&��m:U���
�_�2z��?Ϟ�T�ׄ]�ST�>$�@SF����dW ��بbK}���;����Bi�� ��e��N�J@z/��C��o�Um8���O�`l
ρi�r��-(!�~���r����34�sr�DFM�+�jʯA_^�i<ŮQy
�,�`(��+�y6��B���}�~	�s�\���]��~]�k��_g�g>���7�s��mqMD���X�ˉ����J��n��*N��L�*��\�<��M�>b� �%�AP�=�3����	����;K��fV�r_"I����4����d�.I��f�@
�Z�����U���0O���/ޔޮG�_,���|�f�Ю� �Rң&DF�by�+v��y[BroXz<�kfL���<r-��h��pJfnr��t$7M�=���ˏ4ϥ���-�FsE��,xe����~e3TQ
���O�-W{z��MR�#G��9��2�O��M��=�9�U̫t�jr��)�?���sy~,��C�553s^�b�s\���O��ϴJ�S:�=P��#R�{��ˡ�
���'�~r?�Z�o���P�:�i�m�SذjE�$㴧���Y�_z���CłM0�;n-��3���ι+�T�	�����;cs���U�G��5�G&�.����$[��'h��PQ���j����0����oX�(��Z�N��P1���҈P�y��7�t7��W�����o҆�;�N�2mDy�藺�u�o�x��(ө$��v̛*�X���ƫɤ)>v7�F���y\�M��Q����Q:$~�W����;��,��Э
�cD�����LK��ӫ�����k�g������Z��~��j�랶������̹�ʥ��hh�K�/sv�<<<l�7�[�o.��+�7��.H�_j@���)U7�����3����M8/�v��E����QIʻ{�ԍ�L#�me����
��l�ǄN^������g�MY����P1�EoE�M��ߏ2�B�'C~Jl�������D���{��`����X��"W��R�^�%�y��rϒ] 		A8������y2=P�T��B��=��o�Ӈ%�m�z��"�GH>�D����B�鯏)����,т�vX��H����J�'gI'g=w�Kj�ϟq<1��H�b��X��Xe
���3�a/�X�9;wI,{L�ӻ���%~ �D������ij��V��V�3�+��U������2��X��o��X�i:�G�������*V�R$�'��ݶT����$���W�V'�=]C��XM6e���^�y=.�Hmcb�1�^�i��6�تK2��,�ξ#S��%ک��N�g�PQ	���d��,�O�9�5���od@��,kw$�/c�x�h��KL�:7��,�������;�%��-2�&�35���s}�Z�K�������H)F�fe�c��o���9g:���엞Vx�]�D�
	K�����i�ܯ����>����Y�����/-AtƢ��1����K��@2���4���~�Ġ���"�I+H�d��k�#":��lؒa[aW��g�@���BW��3A(h�a�!����Unc��a�~�/�W�A{��hr=N���O��V0D\BbN}�����]��'ʼ U�������W�B??�=����XXa'�M_��W��9�p��]�&�aI�er�f s�e�Ȍ/��ر?����Utꊴ�eT>A~�W�z��3_,�߱�̮]�����ڤ7��|=̆�w"Zq�S�Q����8�������$��	�i�GH�g�o��,���~�(��{�:mjq1*(]J�4�f��?!���.s*����SO���������^���^�l�BJ'�u0O�݌`t*Q��\��D9�8"��Ҧ�w85>�ב~�B8��#�a����-t�sTl�;T��i���o�GR��)a�=�W!�dƕ��1�6��}�W9E������� .%u�G��;͆�,���w5�{Z�s]XI]A��/IP������
��؟���f&�a��0���qT����B*����lo��̻��>-,��ch� ,���x����@4"bP��GU�~�V��T�L�X��Z]5 44b�!�g�>Kȕ����oF�J�?�;l���*����ϟ5�h��
^��h�N�QLf�)�fon�+CBvy]^�d=U��QT��%;�E�$�g9�]�P}�4��"��~�?��ay�Ġ�)E���vsv)Lo#�R��;�q��]��
?a����R��P-�:�* ;W\�V�x{�N1��;�����=�E�a�յx�I�GO�[Qx'�AddL�)wٟ���lz����ubb��)G&�fv�Χ�Dx�(�Y���I���6�rm������ 2��Cսڊ���t�d���Y�'�9Wo�9v)=�u��0E��!����(<������V�*�\��g�NP.��V��=��j��u/��Uf@�.Ǉo8U�	��U��)�5U�Z���� a�2�6�t����{��6���,m϶D���t]��	Vb�w�oV4��q\�b��w�­s�
�50���oT;�� Ki+�"�S���>=>MY?-'���&�ߨ���#Т�pRR(q�4�l����`����r�i����E����ׅ����Ȁ��H�-� �Rp�K5+%�J1����&^#���Z�C�4�V�$�TTb���Q��D�)Q@'�W���n(=�#J~�hn����)���0��,�R�4-*(�qSP��,׏�$��%�����S�Vﬠ�j��H���	���V��_Q�L�	ڂ��.f�������2�@���$���Q;<hB9��o���iU��Sq0�����8by�ݽ?ՕyR��L��O�YY�}�Qf�k|Z��XӃ���ԟcs'0FX~�,��:.��~�(�� ��3�^io������&i`�0={f3���������҆ Ӂ�n��\ƣ������ۓ:JK-����z�M�ү�I.��.��C��(UP��D���E{�X`��JH��L���R����;W����s"A�)̜���
����[
��bq`������P5 ���=�F�=,�>O���Sv�yO.dP�r�ϖ�-���V�䥌Ӳ�K�ĶD�g)���~)cW$�PΤo�j��b��}�H�D�a�+��!���P�T�S����0J_t#r���K��X'6���^St��Ƭ��u�Ĩ�\��|L0��1[Z����3Z(�Q[�1ſ66&���o ��7�h�l�����O���bH�����HqrD ϲUr�d�҅�8�?�V�8mD^�h�AsP�9rC!��m����B�$)��A�i޸J�l�����Gi$��A_p�
xw�@IãR��3���t�ᮚ99��BZфK�<������*Q$V�����L ���˽}?I�48�Ѕ�l1�A�.z�ځ�DC�!�;���ȅE.���Q �/�,3YO����Ė�QT4E��H5����
x�ݏ �b����=��ۯ:�֥<>��w�I_���M�v��l浸I�I����,�wX�BR�(�tB��,����2z4���04�k���\j�l:��4���f��ݨ���CA�p��'G,_��l�z(�����FZ�x���H8Μ �p�^�q�A��yg�7+���W��pݔY�~�R��Ѱ\j�ł��ۤl�N�Vͳ9E���#���ױ��Ww������}�)$+PCC�}���}+r�š5W,R�G��!^�zdD*��C���#����Y��_�	���W�Ȗߵ6��w�D~�zo`��Μ(��~g���8CA��!��~���������߽(f�����zh��(qj� �L����y�oY'�9M���ҙֵ\�+��jl�,C���k��7�/�hh�:\��\Cx�hE��?��Z���p�A���_< �Jq��`�'[��`�{�6r�쬱�Ƥ�vݬHq�nC*��������8d�����)�X$�h���`�����\�۶@؍�������9�������۪h��j;��UdFc��A��;D�ԃ���){ARKFFa�oI�n7�jc��Wy�dt=`�i��ao��:2������M�(�O�f&�Sepy}�'t3h�B�3w����
�T����
}(bt4eXh�Vzo[4��Y�T�.���S�U�U���(���}M����ۋL~x��R'��dtό���M{�� �,����zf��a�����=�+�1f�w �e;.Z� )5������f`Ⱦ��5�#yĀ{�]�$6��oHQZ��2�Ra5w�*������C��l����̟����������V�<}\��Xt�z��]�K�[-�W֐r�%2A����yt�I,��lb�r'��F*"��7,VŪG�OV�q��ϟ?�}�`T^U��g6�ƍ܃Y��̷��>���BV��G	/��-�.�N?@���)w*M��Y��\��t��x�Plz(�xeee�N����H���G�T��BZ5>�{|U�K��������uml!aÄ������oq���M֣�]'�4��+�n:ZI��s���n77�_꒤k6�_�2�^�ۄ�.���pN��\� 4
�hRq bJf��x���#��'po�"!��PP�IW�����E����Lmț����1�)vJY��'g56�Wgj�B�V
��y�pmd��t_d�^��ή��R|��Ol�=�%	ÊH��+�.k��R�H��[Y��y�m�	����~����'��uU�'�I�æ��N������'�i��8��E�䏨Y���W>��o}��+�����vY�S���0���[�v_���(nŲ!��w�����чָ�G�fA�̨�"ܸ녝��|��8�rb���{U��8��Sg��;��^\BB����݅N$#B�g䒋��c7>��k���`�Js=�6��<ۍ�]��e�6���Qw�)Y�
ܳ��ǫ��ї�Tf�2.���Ļ?�{����d��)�ҒR+s_H�5�.D7?O���Yhv�]2��H�@ccӤΙ�P�Tl�P����Bn�m�\��m=�C����O⢯�4Ax,z\w霗��������]�ۭ����7�M��}?R�،�9�!���jxk-�)�� �;����R0j��<��V�㾨p��HF���&��'��T��aEn��c ���xv����WuMr_L�U��IŨ��F,kͻl�
Ɇ�'��z�W�7z]��:I���mO����:\���6V����u1H�I�lƪ+���:�N�� ȁ�|��1�Bj]�'*�>��j\�8Bӟ	 �|#�Q�T�<k�T�Y�ܣlճX�@nn��".M��%=�
8=��^��vS�A{ŶY:��7����`�!�7C���m�[j�@��kj�~��N\pL?�h���Rb��@ͨ�_��AQ��]�\��
}̾����x��k\A���q;�3W�A�n�E7��C+��r$%�ג��kym��* )��^�m��H��_��|v��.m*�����O��Ms����C�}�.}����э�Qg��h�J,��� �*��E
Ճ�����ī�~M��`�m�]��ͽ��@9�N����,ї]H��\��k���b�홞�>4@��}���B ^� R	B\��AM/a��yo���&�����8��z�*5Ɋ���?N��M0h����4*�n�=-4�� /k }��������8�V�'�����<�`ԏ(�G��]p1��\�����o��mx�7���0�[�����y��>*�� X��8�\X�����u�8L��-^�#�M�tƉm�-��6��/�r�l 6����3�Ѩ�v}�b��χ�Oӡ�A���b�8��˗6�F�}-�����b�B=b�y�h'(6b@Fn^t���g! ����9�@���[R�g�,���,�=�*Þ�.�����(���Y��-U`<�ж��U�<���w�����r�$��OX�"r7��R�J�+�N��JW��E� ��rB�xE� ��,�y�q����<~�����*i�[4��ֶ�N��ӤSVje��oPgI���|������/�S��D2�<�sE����`�&$I�ѱN�p
�*��{7��o㵶(KI��;�F���Ԕzʡ���ۮѱ����ȓ"�ű��0;"o�³V���P�R�[*��D������^���8�����p�,׳O^j2�\�����H4���Uyy_�_���9�_�n���*q�2Tc|�#�D����0��s9�y�;��-��(����d&xz����[w�v�_�@�H�q%���Z��K�PTbJ6�c>ʲ�n�ݑmwD�x/�.��g]Uc6NN�����),�	�>}�\�M?'�-׭=*üp�]o=���ៃ@W@��q�H���,w'���{T�ǌ�#�Ɍ݀�*Q����m8��??"
C��.0* �<lҊ[�U�C�~i�V""�@�7��;5% �j�����[�Ő`���48$��u�ϞZ� MƎ�+$�fXՋ���!�"���&xX��ߋu��vUG�,��&e��g69!a����M/_���loG��r>uyh0L;.���V��5�`��U<9`0�̮�缣�Y�� ��㖱�k�Ei�+y$#2��:,���.��8P�x�q��)�B��� ��]��R���v���Oh����QPMa������(�y~�f���vp���/9;���Oܣ�n��r"���!�_�v��QQQ�s�S�ƶy`ع��,`�ҼQ�d���A��̗�﷎3r����Y�n3�Ӷ�'s@y}L��ܞ���c�n��k�?V����������nybv��7u�����2mzE=O����2�
�
غO��* �K.�_RIF���'wsm�{�@����$������aAb���>y�]]�ٕ��55�<��5���V=G�C����!�����yG�s��wuV�G���"�V[�^�&��)��ipP�J9 uQ��GZjxwϢ�!�L������E,���D���;�R�̬��܀��P6���?%�<����S��b��"5!0U��,�����N���	H�&��r��=J� ����g_�� ���6����K�^{�|�`~p-��a��ݱ �o�Jsw�s�:�[���6'N���[��D��� �xT
���������G}��_ ��֐��X S�H6�@1�4�)��nRB@�zݤ[qf��8�{��V�� d����xH�@'p�=S�9Bk��ެg�sLt��|V�v�{f Ķh��U߲^)�II)�2���L:Z���/dT��}e��,-g�����[5�E�%ZpN������T_�j޼{`37�Q��ٖ�]e�N{�$&C�%:���/$@$�1i�|�7���7��L2 ;�ȠS1�+�?�q<�j�
ѿfBxjN�UNB1Ɏ�R�RX��,�$�S��J �ؾ�e6��3�����L�"�E���4���A�/6��ݙ��z����ڨ�cE��ǲ�;{�N�_Th��tfs�ެt�sj��J��\�|c��k�:/ww.d'.Q�KE�y�C����YT�ST��	��UDĀ�/ت��]=῎N��h<�������?�N��V65��|�C� Y�٠|��:=�iO(�j��ۖRq�c�[f���/������]r���x��v;���q�c����|��E��R=T��yc`�MA�P͸��V3�����f���t<��"S�AY}�}�����%�Q֝C��@�{ԇ��⥦��˾ժ<��ɺ��Y��F��ׇ܏w.��gg�w����:+�r��`s����_�Ps���(��X&��f�|[-(���+P��|��f*SU\�)l��vy^����V������8r���;���H����e�ڂ���?��~�W{��� �7e�y��է�J���]VG�mh��� -k�kU�Vp��-E���a����/k'����`�aG��ڡ;�|���/T:���������Ջ��*K�M�t|<��rSa9��'M�'w��U��`:mm�������L�@r|��X�Ӵ�����V�]�<��������~�;�
G�]d3mސ����:�����������Ś߃;㲙y+�@t�� �ޘ��}m�ՒƬT��_S�N�K_R6LRs��l@�����Tl��~rI�C�抽�{tz��5s���+	@4��3Ѱ�ok@�'�߫��q����^_#_��%%���|����#��Mqh�49%YS�ޙl�o\�N#4�r�16R��kX6�/�9��i�$�:��߁��!��U��s��kI�X��ӲB3WeLo�栣K/L���R
h:�Ra9��j�R��{i��{W}�p2kEP�uH���z}w?�ξ�|�@(�w�I$8���6���|?�1�;���qeyJ��ȩ��x�V@ei�M$���I�g�P�(�v?� �ze��|
7Qv�����\�P���ݷ��*�F��S�(ۭ.ݕ?-m/ੇ� B�6= n�`�V
}�e	K";��ev�B�d��:C�%r>�����z��gG�،K���+:�/2�P��1)���>�$C���fo�^�?ֻPz���km�ܺc��n�uc`/QcH���s;_��;콃�գ�:�0]�*: =�⬉���(�a�ld69���{�Ғ�O�V�D2Z�� r��*�ue�py�xl�ɳ���K-�ZZZ�eR ucOa�'-��[D<;�Q�%
��HM��J�K��{��DM���Ǆ|��F�'t�s�n�Vn��G�{Ƞ�Ty.�'ЋLޓ�,e�����}����mo&����0{�`2˸�t�6�����>�P;��DQ}Y�hk8DLS��M`8\�?�LK��EEI=O�\�vu��E�����)�R�/�~߅�������
�u1}/���J/��\��-�ƪ�c\�wH?���uK,��]�G����a��H��^>�}�4l'7�H�d=,z��e���J�����a�$��?:4�=={ w�X�;6�@�}��L����˚���e�%
�j%j�� 'R���
�<fs�&� +�y2(����.U�x�����M��j�wɻ��j�3D[���I
��UU^�|n㷊fK]���w ���м���%��}��\A���kEP�|�Z�����qL�D��-��+
���ߙ���0.��=�#0 �6�u�o�8��}��̴gƿ�:k9��lKw����0�����ܻ׈�����������8����l��)e%��Ml�'��/��l~W*⯙ɝ_}��ٰ�q~k{���K��bP۸��;�v����L.j]�AC{�/]t��;������{쳘<L�ӊ�+�
���^_����������`�͎4�j^�B=6j����_�QsA�Id��|���CW���y�aY����Spq���Иk��ov޳l4ί���sK8Wa�Kz��䇒�����Mu����'��l�]��E�8�Gr�Ϥ����[�?�#��F���Y]���'ONa&+��?��f���@vp��C�o��a�{�R�@���� ���:���ߩ��U�v�ڪ�b���~p�P�3�k��Xߡ��0�Yuf�#��� λ��~7=B�K����MXz�v��DDҗ���ȱ&+�R�!�����GVz~�_C��-�l������Y���:ԩrŨ�������*�����zsE����W�^�1ъ]%������A9��g_�m��Ǔ�,��i�s[��&�f?�	�}�X�<��G�c�AZ�t>ʇy�hD�N����g�	#���_�� ��:6�(B~�,���,T�4��G�k�_��	����p1ǭQ��;6fG V�3N������ �I�!*8�\�EM��P�p�\�E�u�����'U�K��e�e<MvN�rkj�F�(��R{1d�_`/_���I���݀�X2�$��5�hl�x�ٞ��g����.���ｸ�T�m�K�JJH���O�(�~
���7&F�8(ތ�%�%	���[�����6g�R��E�A���vJ5��vZ������`2�S,�b9��A۠sS�pm"V	�!!����`
Ŏ���^�I�%�7�D��=���пaq�������hr�5��{H*���'6�L3�� ������Lا�'K�,IsOծ���\s�H�V�" �=����h��������m~�v��9ӿ~=�/;$�*((Xn)FI��ҭ�x.#'#
��<f>L>�߼F{�+�}4�d%���sk�]�3B_uf������D������`7�[���4�M��,#bIf�T׵K��4��L}�����z�ڇ�S���mط ���x��X�߯RJ\&���X�1�7�a^hQ�z(�m!�s`��Io�Q
�SG������N1�yL'�����������Z����x��i���]�+��&*c�|�ޕ�R��u/K"T*���� ����\D )��T�qq}xTHe+Z�fft4�u��Zz�%�Ӡ����B��Dq|VV������I�u|EH���2�7nC�  ��R$\�:*S䃅��R�&�q�����Z]��Lޱӛ���Vw�P�d&�2�s��qq/�]�g����,��N�%�lG����}A�uߐS��%��8y;�xf��4���ek���u�HNh�u�V٫�s	 �S"�����E��1������u3zwP�[�e�C�^H�ʨS(�^)�ɚ���B�<%[Ey.�^��H������y��{<�	�t�~��
��'2ţ-�>V�A6����ם�HO�8Y�z�οH����)"�"#��H)�!�dl�`@����̵x:}�p2G(��M�<�h����{�E=�������+��U���[�>�V��+������T1yL����[�_^���GL3����HG}�L�Z����w42�Y 	$��Ksq�x�?�g1��ͬ,3*D��K��qܨ���]/�En���ڢ�V(w��U=��`s77���-�Wk�	�� ƒ����q�Qr<���Ehf"�9���c4���Ā�/����=�į2P�6�ߣ�`�6�!��� f� �-���H���{�/��W������ ph��ņ��ր2��־U�t�Ɗ��Z7G��}3V$3��@h��X|���.m��Nͦr�\�Q�߰�X�a4-]1�JYn5���sc��<��6����d�]�ps��K�������qΧn1M/@�b�%K�pX<�'zuv��xWe��[�<�~AJq$��Y,����q�|���.���/��΂��:b�7�����'J��H���i���U#�"����$=6�z�+Nϝ!��F��,>CGS�  g�׆|�K<<�.c�'c9#�>N ��>~#�+�2��T��Wۃ;�����������c�-������L;��%��~o~������j�x���m��h0�	I,�Z,d��"����/�s�g�`�z��$�=�YqO:|����fi��>F��Ü�IH3�D��7��߾ԃ��9�>��e{x�������/8~2����w�c[[[���R0�����<ɨ��3o%����X()E�?<X����ky���)W�D�1�iu\�/yoec:�A�x�6��9�*��r�Y��n��s��]�,>�)�_i�i�V1�W�Wy�g�����m&4�:���8,"wja$Wz�Kw~�ݨE�N)��f�ԅ��'k'�)��&4�[wnM{#���HYYY�&�A��`���C�T�*6Q�7�˰s��UO�ݎ�'�Z���i�������3���E����䛣����V�VwHb��Yq��NWw��3�kw+����^�.��{���M����Y�ҟ���g�#=l]�<���j����7[�,��ق��+��||� �5MVv���:t@��^1W����3~U�Cb��ùyd�S��Q�L��p���� L�+��uX7t;S�54�n��7?V]�٨�P"�#yo���CuW��#IC�	�@�}�UP��i��㕡^~8�k�2�0���L�ǚ��-�S��SУ�F���7o�$;QE�`0y'j��f0�j�<���iy�I�C&��z�*�v0�G�c/����޸��5���{o�[i���=�,�����.D������$< ~��YH�� #c�/�-U��F��g�Ve��*v�6�Q�b�R� �D�&44�d�Hq{��|`bWY�Ƽu�����麬f�u��*������׊%{�vEK�h�!!�1�+�0㽹;>�����Z�d!��-�p�T��U+K�2Sre�`�	r��!⥣Akt��6�S]�_`��3GϞ��MPDyZ2
H���ӛ��:6�fI��q��0���a���nYG�"�g��3����H{Z���d�� w>��%9l��ؘ�/��j��۶�ŀ|o�S����i�@�������^��Fi79.*�n@{��O�&h<x:R�>a ����s_遮(�M�.YC%9�35f5����&�8v��I�&�5�����
��1��JlHr%Q��]�-��g_��7U.���p)�W�FX�h�X�����70Rc`��#=U��Ν@����I����lvwy�J��2g�Y.�,I]�9��k4�_B�~��ܳ��8[�����uZ��Eםq�����"�tN+�0�����rZ�ڦ&���\P�J��������a 5��u^~~~�©�ü7�<Z�/�BA�B�J���+�u~j����𻫱� �)	���. 5c��(�PE���O���]�'�+�GIXI[����y�7:TK�lڵ�Z8ssED4ʾ=�,��v ʄ�����_+�},)ah`]����F����6��<�)���U͓@[p���m:�sE���ad6�$�6�"�c?!�����-.E�
�:|
[��~�W����u�'��mx�q��l�Y�{-鴸���R�& 1�1��<���y�\2��5�,��#��XUG$�
d�ԋS--�������� ��j(�yH�踘� �_�����SD�_]R��K���g�R��J쯏��4����t6���W�kL{�cx��#a�\��QU@��@ұ�ܡ1KKK�n��s�+%�~��5�%V��pP�d��t�,S4�pV��*`�1 ѪJ=$�UG���ه��Y�g(~�LA�"z�z�;���>-j�i\ �����f�%��.�����^���Oɧ�:�^y��+��m�d:o�=�F� q@�iT�A�t�]A�;ㅻ���f�F� 2qہ]�Fu��ڹ�_���}mt����ݜZO�]���["d$gՕ��W�G�;�O~��Ԛ����ޔ��d�`���Zwl|�㸩�c�'pۡV3Ț0��<��[�,l;���u�<���׷��\\�/�ч��YE� �Zl�~��>�� ��w�!�O� �A���X��eIv�nbC��߬zs`á� U�3����\Q��4�@ռ���LC��.����BM-�������aQv]����tHw	����Hw��
Hwww7HJHw�twww� C|�p?���k8&��{�y������Sꟶ�{���ٍ '�BkN�a������H���r�� �-����q
�;T��;]<v�YosV'��H*[�T���~��㖗���S�(�w5L��l:�12Z�Z���!�{U`妳���m�L�����)�|$�Z����;.�%��_�]Cɣ�ѽ'�u%��T~�8�F*?<'R"�l94�g}�6�z����KC�����C��F��)���Ք�&��Ĭouggg�`:`���KH�(,0�d`�(�%B���l��Ouj,P�t��O�p��I"I��t=��&��%���5�;ɓ���d�h4yy���:7 uƓ�*b�o?�lA$a�[	,+^R\\�pbAF������ɔ8�'Hӷ�l1�g����@^����-�:�i�O����0�d[��LЛB*_����$`)ڠ�9(gv�7��h��Q�󋋁q�\�N�BN�l����-}�a��Fc�v��6�����Gá$�ov1ֵ n�/�Ŏ�'�s�hpە~�=`a�����°�zF4%� �.�Ŕ�ohHn�u (��7!�Ǭ�l��o?���L7v�M~��O�8�/�&�G}{��; �$�R���HH�����za��ڑ>��2�˟wڷ���B��Y���Cq�G�q��m�,J)���a�J�$�ӆ�%���7�/���D
>q��o���.R��<��L�����a��>Y�݄jkwP
��vDr�XZ�J7f��_�� �-�Bg�֣Y��T���s���ǐ�<�˕��R�B���o�>~*$Hu$�O������lW�I!GfC,]��ڨ�3����SR
�}����O�XƉ���<o苞Q����Kk�t�5�Te�G�g���O:�j�`�%0�Y1��m���9'f�Nk8�L���L�Ɯܲ)��Oh/!�C'��л�w�6�;$ЇR�漝9��I�{��;[�1Y���w�F�+Ju�'���x5Co�/�v#�Ūm8CPpz�B���`�91�!{���.o轝���T�ҁk'����k�� #�>���' !)n�2D5�:�훝U�� �-�ϻ�m �77o/nF
Z�_� �b08�yK'�¼��U��fľ�Ӣ�k��E	�)������Rmv)�������n�c9-ӷ��Y_�7����U�����v����c�Z�m��0��"PRR|�⹣�x`��#�9�]�����������6`�Ś5�u�u����<?Ȟ^�O�Fɯy�z�JF�%��/a�9/v�#���
��Ql�pWX�S�&�h���W������?_�?�B�-^���GY)�C.$O�j��31�e v�-�I2xVV��]WQm�>m'��˳'�w����IHH�;3�S�����J+�a����s{��I��hSa�юgs���ES�f=�ڽoOZ�?�+ 0�lcmX��4�ݽs��%���ϧ���A���7tVm��,�Ȓ}OCW��UG4�.�&J��N��-�����	�����{�����/sP�u��-u{����j����\���o��_��4UZ�U�Q?�qb"���[�*d��ɷz17�"z�k�]n��-��v���x��4��Ԓ������1u�2j&g�wk��q��<Ek�⭧��m�#g�+Ӛ׼���*C9�L^:���A*j�Ƭ����zs��!��2����Z�J��B[��)iIGH^�Q�o?]��\��F{�B(��F2�u�}_LS=Kq4)yF��-�H��Tp��x�G&���J.����褼~�u�E���y�V �w'x��.�ª�W�hzAI+۴>z�D����b���l�H�"�f�	A�c5�%�s�����֤,�ڸĠ?,%��9����7��w953�m��'Κ�2�?"�S�� �7j���{^�L
����x����u9v[��lB���Z�B�[�<K3|�*O},�����qp�=�'�r���S�p� �����z��*\�Ɗ�E]��1=Q=/2?�XIL����T8Zկ�PO*��K���{q���N��)�/;�a��b��9�&� �D�ϥ�j��9T��Ɠ�����x��g�\��7����û�\S�S%��$�
e�y�>\�N��B���z��8�d͗��U�Bϰ�02�5'W��[@���=iih����343.{�(�C�;�C�[K99'g+q�蚘7��2��DG�b�޾(T�'����4�L�O\H��O�m|x��dz�_?�	�Ã颃��(')��|�\�9{��5�5P��'���d2W��z�G">(66�kd<�����]m���z\cv�Ms<{��~�J���.T��"�~��a���G\C��-�QùU�H5�qe"��T�u9�;��!4*�	�,��nϧf�o�����P���G%���1_A6¹�3,T�_��?�;B�tbSEǆs������Z.
���*�dB�դ��#��u�k�T���G3��S�d̥�� ���=�\���~��lKւcGπ��L屝r��qH�Z�r���vy~z4�S6`Ԫ�?�JR���3F�%`U<�Z`a����7ۃ����X	��!!>+�F�zP'
j�K�S�Cc!��M�v+�<H. ʸ�8^j�Vw�����iC��*��"�l�J���:99)���y�^i7�=�c�l��:{�j�*�W=ͬ{?���d�͗�B���iMP�:	���yG]G����;����uE�E�[#��3?� �n���L�2��%<�<-�Mq��X2�=�id�[��ч�iE�1xV�%n%\yуٲ��l1= �� ���l�=T��J���؝�.G�?����P;-7��3�*N�����m	7�C����-�tlT�u� �O�Ym�imk���"Lƒ�!v�S<��n%$4T)�ש�������9<ֱ;88PPҹ�H%0�U���0�Foa�\;0�pE��Y���~e�as4�KG��z�p������R�6�0��(Գ&�#�fmM�v?�d3���}h��	z#�{��<ȣ��Ǭ�9�%������9K�B���k��٤�@nEo��-J�
I.Rh?G����pZ,���RUz >;+7j����,"��DUޣ!�z�0��Ѓ&4v�7}:���Y.�(�IU H��*+�*kC��ƄPd���»|���$H���$BXX�na����U�xi��	��;��Ϗ�3��Ŭ,�2��Eh��ݴ
茜��s~|m�^�mh��Ȼ���b3������mDhR��l��Bk_ppp��!���	u��*�$$޽Fx8��G�$..Yi���CFC�y���|A����Z�ƣ"5�x�q�o�m�bǦ�g�Y8�W���+��.��XK���[[U'�YL� �<�d�?��z���% ���_9;];=�T̕�>�@�ࠉ��_r^E�YR�m@�1q�֯ߺKm/�櫖--/[ߞ��}�������rvq�b�/?v|�з���=���N3��:��[��k���wOK!{�����>[q����9h����5�|���w{0Q���Ze+����Fx�J�����zm��oPP5��`H���UƁJa��{J�'E�|�^~L9� x�)�xce7t'�=�!�⹋3�d嫲�G���������o����!QNHqa%[�i�G�?X#�yj,��<<<����S�͖�i�i�����)ր��%��57ߑ+uv^�)&���b��@L	���j��X���UxW�^�u/����e<㉿����JO���k�ݠ d�e^�r��Z-A���
T����ndd��w��t����꨾B˸��!�,�-��6���������7h�1�9��ş�������1�K�(���|���c��<<���V���"��*����2������6U6�B�ݍmjVV���62�����v։zmK���ٍM@l��sQ��i��`-;�[�P����ʢ��/�`-���g���S��A�U=x�������]E���>2	��2S��������յ��I��Wsi�րW���t��t/�>m�)3�b�F,���F�ŀ�(O-���vkE褂���d��h�p���b%�ͷOv�Zy+�o���f@���k�r�_81Z��P��a"�zɊ ���zh\�RH�����>�\U�I`�W��(�����g^�q]r,����ׇ�ԟ��994��A����H��{ӻ�b,�F�W�볘��hE��qp�b��132�{yx���m�F�:1?��ٲr%%�5�m �ؽ�ٺz��a�1�(�3�v����)
��8e���f��X��������1��l0�p����9�4�}�삣�gW=P(�#�}���P~V��b�J�r.s&Y�8$��Q��8�)��B�V�[-Ԍ`��t�oq�;���1�?�W��k�S�
и��o��r��[��l�^�B���olZv`����_�L$�;2��2w�����JS�W;�Ƚ�{�-z|P�7����E��ؤ������u;��=[�}U~~Z�^~����R�%x�����ʩ���w�a�e�8峧�rp��쮔�${��"��`���®�#��z������\�OŇ9nK+>�Z��q��͗��be`ˌ ��b�Ki�M8��獕lv�.;�}c�A�+\|���Ǒ�Yȩ�Zb��{�?��Qs���4G�@
�~k8j�pvH�*��bH�&nt𱀳������	�5� 5~��.}-�����{�J	ܡ��ߢ��T����KJ��N;�tӍ�⸓]lez�۞�.�g�Z<ɯz����H.�?-!�8�m�_��S/I��g�\�t^]�'~��N�/��#/��7N�T��Ao-��P\�_ÛR-Dh+=������l�7��d��Ԃɳ��O�V�Ƥ�ԟ�f�1��BYګ�����z"�f9<t*	P�����^:L�m���+���E�M�$dTT�8�����҉�n���h���͚���W��x"�����=��x<���;����pH��ߪ ����:w0���v��u�H:������yH(�c'�2'jm?��L�J�����0͙������DNVBԆ��P�4��`Ї����y�e*�R����F$�I��oz��؛s����|������p��\��!lg�}[��b���ht�1�9��#�]r�[������4�\���;�nhPWӻ|�Z�>�吰��Ҽ�}�Q�.�:ʨx9�fr�������J�"�����(��,Q�a�����6�nv�T�'"���ʐ�ۛL�1ł���f-�$�=�*��uYTT��Ϻ��L����Ocb�R����I��6R��ky�B�Dri~4E���j�ҙK�c�+{,�̓?�Qo�ۛ�Ð�۟+�⒒>S��+D�DU��?�N�6�	v�ҭ5andw�XP�Y,�p�L�c���cPQ��,}�GƵ���R� ?u��ǩ�垬�����lJ%���^�-e��Jv�R�h�?>��ʓ�y����dY�y����5=}K̊���]�#��b���E��%����W""x��Z;:�0(��8�4x�s��#�2�J�O$1��Q�'���ߐ���p�[}~fbݢ�������#�yX��2d�t����K.-���Իr&SV�Cn���M�n2���a�p��`�i4U�g^���N,`	��x記�/I��4Rl-��Ԩ�C/!o'�@W�E��E��D3C���u�N�#}D�4�28m��'���X��[����2E\����[�ä���GKu�֖����;M��e���o�О-[o.�p�����z�G�R���ʈLeTmE����7��K5'=i��C\g�I�=:F�4��]�
��~l�u���}I&�]X�g΂����3�-c���,�
�ǧ�3��r|�I���]����;��6�7�I~�9�"�t�x��V-s���6-H/͖����'���my9�Zj��< �g�HQ�X�cg���5���X���v�A���&_Z�8�������l7�B����D�J�o��{�s~ef�n� KC��Ugg��B�-���K��������/�@l�� �Jbsp��Y���f}��=�֕�M���=�l����0��r�qL'ވ�¡���s��Ʌ)�a���p�=TX��q_~�r$_���$�wJ��q�$=��o���ϟ,����RV�u��)���e�_Αk�&�y$dc ��޴<Σ<2��O�G]'kf���mn�l�xӓ����~��j}f�^p[.��)�4�����'�X�s�]���ME���bK,Y�k�v/����H��̩Zׁ�k�z;�a3|2��ko��"ξ�3\�N�	�2���-~�U����������JH�=��"��'�kΛBx���,cG �h�Ҩ�S��NO��|~.��첷�kۼ����{�FCXS�$�U���?J��#;�Ӯaҗ�,������b��>�ncU$5�!��բE���>�xV������b�ࢌ���H^��KoA��o+�S7��_h�͇�s���5yUo��x��P�XRW�6�e�};	38��jғ�e$kJ�r.,i+�)"�ۢ��]�:n�[+N���z��F3G��nk�xh��h4j}��l��H ;��9Eq�n_�������/�t_nYSf)%i?�׻������`0}ɩ ���ʟ6^gu���uW��P��٫a�����x6~�V�b���V��)�����*0��ސ����>?�ծW'��<rn��C�8�5��`�e���4@��ω4D��g�v,��1���	.PP^Bt�G�Y�hq�
-�
a��}�Q�м0�崤Q�ݷؚ�ĆV/WV+���qp]^�λ�^���W/��ѭ�>6A�rY�S�TP!��,Ϳ�9��":skt����!��jd��ģ��i���>����~�Z��h��4-�˗>@潎[c2�s�Yݼvq�L"�}T~��iN���3(50Pn��2����i��/�BC�`�b�tX��ruz+/��|��Bf�{��P��H�`�	6;,��ZO��N��Qdg�s�`���]ye�4W��J���)X��Z��m�Вq��fT	�z5dԞ��d�l�?��h4u�&zu�L<ي��\��"�d ~�ݦ���u.�*#��y��FvOO1��������;� UN�{G�	�c�߸���?&�:B~H?��~U�?Dsr��Z��##[?NY4�����t��v>�g�1U�I�y��z��<s��!���3���֟n)O��S�����qZ^�{��"G<���

��Q�s�5��'k�!G��V��������cD��-�b,Za��f��#O�s���I�]�����X������]��
��=���Ǆ^��`����&6�E���1�=(r�����Q��\�{$�5��Y�acm�����n�㢯��;��[:>���Z������{W9Cn)Zg�h�9ɗ0���f�|hnn1m����}ueǝv�.W�kؤm��y}M ә�eyrU��H�#��@�'k��P���L`P=8F$󋌌<ڴ��vd���Nk\��O5I���j�Xl[�Agd2�'�=;�"��V�o͗��.*G{��<�!��}�z*m�R��R�΄����[��1�����K�:e���b�N���}e-�?��P�����ذJ�~�N��q���� ��%^�ك�WM�_Hm��F(��iN�i���8Qi ����SL��̀� �[���`�p��h���v�9����tA��f(�/�q��&wN�������o�+��)󕸥�QM%���?�&Y5va\�Z���HJj���j������,/b�Ծw$sg��5_E�5\�%�wI���2G�E��Y�* /�&Zee�l'�[��L5������}���/�Ip-}��r{#�l�g�o:ڌ$�� �,�z�߳�lo��v�$$��pA��sc�k.M<����K�u��s�`�E��O�9��߿�J��{Nb���`��#P��)m�9������EK��0dc	h�*?�%��)L��=��$M�
���=��I#J�S�����z���[^rwu��Q1:��[��|�z���H�
�v������{��\��F)�zp�zz�c��3���8��M���uR�[�M�K�lK���Q<��@얉K0Q�Aּ=��)�<CP��'��w��gm���3�M��m|��)K�-mu�y9����Ⅹ1�u��+���'GX[[۪M�ņ��#i�u�6K��G�<����שA�̡��O8��H\A��;��	!�4Eʤ�i�����u��c�1euu��מv�D6��|z��;�7�Dd�`�^Y�����tX[���ܥ��fNH��n�|�q�򇋀a�WT$Kfrxˇu����x�]��������5�B���z$������N䭛g�1��_�ܟ��~`�}1Qj�p�VugQ�n���kq�� �1[x-��qA�� ��Tj��.X��l�D[ꯪY�,�'d�ڄA���ϙ��i�s��Ζ�ܫ�����>);���.� �N剓��J��چ/E���oS]�������3d��|E.�f8�-���3<��?�����r�,]^Z���;�)�jE$,�'�?���>���,ܐ}BAGA�Y���u����B��G����H@ %�����p�Ҩ�UCd�W��Ft��)?�w	ʲ���pM�q���|]݌PfO�}��K|m�Ŕ��S���E��s�Ǜ�@!�g޺��7&fS�n�3׻��T/��坭�ndm����$)Wu��I����9t�{�h.���R��F�(^mBie���C2���k���a�麦2����챆0}�����0g��L�+�c���Pb�W��nՊz+AC9�B���|��	9���bc�S�r�.�Z�|x3�7v�G+���	ID�s����Z�Y&78�L�p~sѺg���	��ew���a�.�o��5�G���6�l;ԅ�|/�E���9��9�`���ŝ��)xڒ���S^:���X$$a���Ca_��$��?u�\1A-�P)����a剨ϊ]��Oq#�M܎��LC�Ie�[a?���J��oGU���cK+U�ś+6��4$��6��>���������l�ЇJd��AF��Ōi?-��5����_��^&��=Pp!��'/��i����9�:��p2�����ELUu>10��=�^�Lo|�7�� T��6��u��(lk��؇�cʣy��$�(&��#*x��C;\��g���w[Wo�$�g�z� ��jX��'��� h=�c�-����t���#ɏ��K�?!f��X�:���j���sm��kág��xa� ���zZoB�H���bP�	�O�UP�5X-fl��-FVD���/��Vr�N�6Ҝ;n��!�F�i���ͺLm�z��g�-��������x$�i��T]����n�$xO�c��h���nY^�����\�� ��� �5}E��!�X��d���;��p��C�������5���r�ȃ5��)o�o�^_'
VGƢ�~���	,�2w�Oݞ��s��Nj�A�A�����^�G������� '�'�w����e�
����Ina���%�.��y�mb�z�JA}��a5�R�u�D�92�5z�-�9�q�����#!����oJ�5s��Y.D�;�x=]�~qrZ�5�2�Fp������+�s����o���Ƙ�Q"S��%���x�<Q�8@l��M��Dk�7�/�ң������&�	��^褩�+�@O(��320P�:r08Z�����_�i�J�whe��eMY�:���6w�9#�+	�깳U���Ixl�J%�+��)�L�n�N��Ŧu�j=� ���M�� ���Z�x]�-�y~4 �臫�do�pF~�{$�;��Dqot���[�99΄k��&x~d7n%o�����l'؅�8�Q�t�E<B��v�PC4<<]J����J-����>!$��ˤYmuw��1�W\���\'TMLvw���4qo����{��h�5��t�#�]�7p���wt�hL�7�X�PV�C~e7EV0���s(��Q3:�����;8o�w�L�)�������$������_PJ�`b	�,!����Pm�&O��Ee�_Z�J��h�0<E@��KA�Bw\����{Eı'���O��`s�k�j�C����LJ���9�-��$�t�t^/��S�}��W�̶��ͼ4�3�ӛ�Д�G�t�qb�s[��=�w��j�_�_�s��g�����f����ǋ�5�a������:�S�u������v����d�\
�5��զ�&�Ϳ�!40��{-i� �|}��I�=�nK܋|)�����O�^Ueꎎ3eb��^Z�+D�ǂ/����/,G�j��þ�Qԧ����'c�W���N��yf>*)�.���T��j�M���WȀ��x��y��j���xB�#)I?K}n��v�,��#Y���Q麗K)ɭd`ףł�#D5�...2EZ\�;v�fӅ�����JLRMf2���Q�[�6'h��[S�U�f~7�`�����p��g@��EaP%��F60����ݾ���w��?�H��V��w����bI=~��e�ӧ���&A�5o`�E���+��Es�T�IpZ�dQw������2m�>,ҧ����+gd���bffqֈA�-Jt��� /~CH�o�'�[��_2�7�m�_~�
���r�̳Ά�����p�~\�Ȧ��
?��o6��zWiC<�$����B<2�	� '��8%���4�w�����oOJ��5UY��u)�r�g��~ۍ�=
~A""�݀R�w���^�ޫ=����Y�򣍕�M;%�@�Ċ���ԆC�๐�!3�hQ>��C���5ָ�����f��T����l�Nn��]��a"w�O�t�)XM�z�'5X(h�ޜ���<8ҵ�M���S�D�[����_;6���T*2�����2[��5:D$>թã��|�ws��7A�� ���!A���(:�3���?rKR�0�56���e�('酚$��n����gP@�{�g����o�|ΞU�`�x> Z��̹R��##��_\s�ZVjֆ}�j���ł4�
�T���=-���Ѓ�kO��F��G�U����DBM5T�ﳟ�>qI�`qG��7�)7�F.��벻x������m��rK��[�;>u|ԇ�p{�]����������`�����p{O����-���������:��~~�����@�!��6a:�C��S��L�U���#���g�A������F�>�n\ͭD�� -=+�K�$�Kn��
�K��F�x6�@ RA�H�Sʓ�+��*�ou�\��KTt�-��i~�w�Hѫ�R-�c&j�� ��}��&5�-�/�w�/��ԬV��"A��U�#�������/����D损:��RB�V?����)<ꡠ���k�ʊ6ax��!L��G3��t���;�^��}q<���`�ɂ�����Ű���U��FZ���I/���)�9{vj�z�{H˟h���a|���^.H�s7�H"Ӳsw�ڹ��Q�%�E��G���\Y�����*^0D���#' Q�30Xm%m.�t�� ���xL���IE��gK�_�?č��m��e-�M<;�;���4OV���s�j�v�a$v	;��k�v��N���JbFr��z���s���?��&��YM�����㼬�>a��p���b�����l�{��L�T>��G�2J��7]�	@�܉.��irCmB""'�E9����kK+����~�z�3Ӓh�?}D�詷8.�Z��2�1/``ܹ$��o[��|���r�=����6�axHT���?��Ԛ
�������or��[zg������zOx:��$�f��P1���ŝ↤d�!Cj�1+b|����b냲:ͩ��K.��Ͼe[薒D����,$���˖�C�d�|t��"ý�l$XoB�"b{�f�sЕ�e�߯�:bw0��L#�0��\5lX���F�$_>����I+&k��'V�HU�_=b�tjU*����3'b4�?<4Wg�Fu�|~��%*F�L�g�zGK+��ZR{�5;R�2�syX1c��*-/��	Ǖ��Bo�%��/߹�^�`9�ظ��X��b�HW���4�x����$^@H�'��W,M���;�Kn�c�W���5����V�S� ����Pi�N������lK�.(��[��	m�Ih�y��v�hIG�&��@2JΌш>���q>�%+ �C�/�z�}�!�xA(�d��t�������~E���������VMQ=��FJ����T��0mX붕&U݁�=j�M.	���v�J�������ٟ�B&o^Q������Ҽ���sfu_&��^��ӛ)�&���A���?pG�#V�&��0��Nlo����)>tuM50������6�.��B������_�M5<�w�� 7������%���wA�����E����/�Q����2������rRy^�VA��[ٟ#�	|�KАU��#�`M�������Z"��G��m�J姧�dh��j��_����^{�B�A��ǚ�'&Fa�$��-��[���?��h�-I�݀��3��e�*��yXC�C�m�Y̱}%������}�o:��ጴ>�c9��_|�Q�"v�ₖ�?����T��@�=کO��G"΍V2�hl�Qh`^��%�fLTu�����³�#���N�k��+
����e�e�web��d�	AX<���̑=��\�o����!?��d�vE�zB����J�����q�ך�]rC�/N} �2� Ȟ���2��5�h�x77p�[��;���»���� �k����uz�&��W�?:�$<��5�~�_1����@>gxI�S'.}x���[R�o,�^t�:'G�^u���'d��#_,�y�E��0Z.C��P��5 Po!�t�A���X�<�J8sC��m�֠�����Ԗ&������KvA�LL��ݝw���*A���}M��p?~���'5� �K��Mj�X�g��љN�]����2٤	r���F]x��.�w������uW{�/�����S<С*Z:�8���T���3�Xr�@v4��+�����c��RsuV���-�n��}T�x��T�d�ťG��5���nhS�g�c�z�*p����w'Ѿq�-%�����|Dp��r������&eK�.�H�з�h��ǖ�������==}ӹ���������촯( ���5t���'��{�~�l�[#���۔w.5}ط�i0�ɢ���R�sKX)�:mo�����\o��]��Ԓn��$��0<�<9�|� sRӉWP �*����\2!�����&���0�l{s��o.Չ��\/b��词�g�^9���~E��v�		��s���SVE���Zgq��{��Re�*�D,q\�s�+���)�f���Q��$V���&��e�� #%S��8R�Gˢ�f���:|�ѝP1}xY�g�w�"0j����:4�8�{��;�`w��+ݏ�y�@�l�o]]�٦�����W%�����ͩR�!Q������*.�tdA9\�MQ�`|Z�XĴK�lY[f��*<�zy���ްg��g���F�zT��k^٤�w�VǺ>c�Ӎ-���޾|�ӭnh����ל�׳����U�*7����v�fJ?c��\y�ϬJ3�V�w�c�]�g��P{@���e�ѧ[ev�;OR������C��og���P||����A6���Q�V��KΓ�g��z>F֜�3р�t�->��2;9}w����D}��/�3��"�H���`=��!]kڲ���~ea'��g�a��3%���X�!�ޯߣ����v�����5v>�\���]ivsg�.�+(��}D8�u���� �Ɛ�(Ƚ�������h��*^,$��K�fr�#&ʇ�)� �>c��8�?t3�V�TcM�?̡���i�k@ε�@	����K�����%Cs�D|��� �W��EkZ5����n����cT��D�.$L�� �[�)�Y�L�F3�Ocbb��)���~��h�ٟQ���?(Ux5��j����Uz�Mؠ���;
����s�<��5U���;�:���4�n�{��嚒����-nN��״Ǽ�T,:_�V��5�-^Y�1	��2��,,l�o�� GD%h��ݻ`O�z��N'׳�w8�'��휂�B+�+�֙�2�hu��(��SH�>����7���Ͳ��D�ij<�X���gfYZ����Rc�_�mk���<?����x�����ZNm7O�L�Ϩ=Z���L�.(m�X^�z��2��Fa�NI@� �\R�g��Ö��"�Sǚ�~}���?1ó0Ȭ[�T��(v��L�n��h�|�.����G�՚��K�o�9��m�<��΃�X�U,��&o�9t����	�)ٮ�̕�U_�h�<�h��U��!ߦ�6*�a��3lm2��� Lg^�-d@�7�I)Q"�P����I��A@	�R����y'�]�l���)u�}����,	A�=��<�u\��r�70U�:ê��aT/�i�y��|D}J���ϛcj�����Ϛ!ΡE�.-:���.�V�S�o��5f���ޓ7n��pX�5�ί:�4 UR)�jC�a�����inNE�ן�zK��w��������Eo������0}m���^�̂đ=ܞQ�� ��Of�Άƾi ��psw3 ���"'
���kRA�����~���r�g�������q��g󾏈e��F$��/��\�q2��Z*�e
�ڭ��l'�����}��³��+�O��Dի/'Iw566�Ή.�X�%%�&m����NIAq��8�[/��k��޶x�,��q��Кć���f����c;�k�)C���0�Vr���$q��� ߜ�C��]���7E�H�X����ަؼ>2�i���Oc����y� hOW��� |]7�R�6lB�������M��<lw���\�d�r���k��w�i��$E�o	h^N�F,�BP�`kn��R?A9$/��aţ�	�	���+H�� ys`A�x��􎶱t�ü?���'�07�(�Fdɲ 7s�3�aR��;�L>�u��a-���r�[��'0c�죱��/F�d�xL4��SН�����mg�H��v��bQ������s�n��$�id5Ψ��"P�۷�f�Dh��!��*�w�Ep��p����(*5/w��+��ę�9n+��嗮���p!A�Z�{�>n\G�݀V�mnR/�g�\�L��#�]�mx���59��»�|�@�w��pl��i?�+����#���T�V�s���QBC)Vh;�<��s^�?g�af�VW8�����?M%OF���FP����l��:L�&5�P' 6_������4�
k�B=$X�Dse���o���6?����-��ٴ���W�>�����}���	���GVT�m�����j�@ɒѣ�~�P�p4�7�=�;$*�O�F��pW)ee��zk�LV�S$l���X��U��A��|��h�V�R�ʆAh���6w�ׅj�^/���������q�ͱ��zp��{��\8{�zVr�����h|��9=m��ѲO�����R����LZ�?�/����'�
O�[�E��d`�hׂ�9�X�ě���񲽷��(3t�뮌"1Ԏ�>���@�'�38z�Ь��<c��H"���Fd��Ӏq�����j���J�>\X
���|�O�M���Z���zW�`�6?�Cn�Q?FX�'���&H���)��/[�
}n X��@����'��Tv��
AhcҦZt�r_�>�����r��)X��%a�a �+�ڕ����f����k�P�HWН��;�!$*a� �0�����������'v�$H�� �?GB]3�&��h2������!��]������O��\��Mr�k�Ð��5�8{��_X��yr�K�u(�u*2�6�Z�B7ֹw�+o�����nf�ؕ���0��y�d�ա b���q�d%m�� ��
3�ᩉ;9��qm�͒ŀ�j"^%H��eYN������%Pv�~���<��-�rl�IW>�K��e�:Ȇߠ��V����F�LO��� �ڙO��[����˺����ߘz'�|/�⼏�?m�TZ$V�>d��M9���O�z�3g��W	���>�X+��,-d��11�5���[A_��/6V��5V���k���6��=ڴÝ�+z�	Q~��Q��H�O\n��ejb�ƳC?��Ŗ�=����k���4܏���5�����ZJm����[ѳ��t��t�2.W��nP؈���ў��#Q_l'z8��O��N_C%z��ۑ3��\e[�،d���E+�vw����ޒ+/�����$����aΓi�Қ��|�[8{��Β�=���"g�N��mC��GIۇ���N�����wN���f���<��]i7@�н��WA}��<��}����8�&�������)����i��Q�V���ֶ��}��$~NB
r.� #��Uz&P%pn�A}P�<��J��=�������si�0�2�����7����/�K�]7��٭Hy�g3WU���h�v�ؘ�*�dz��3��x��j'�H�d[�bW]�vw�{\�X̭yP��G�|R���xv���c)j�e����ʸ���� �-�!H7R�R�*���%��%9t�4H#�0t�P��x�}��������묭��,
�iŭ�$����92̲�j�N�~6��:�4�Y�Huoy�an6�Y]�������f�T� ֆ�N�H�O����n]�Pк�x�&�Xz�$e4(7��ç+�~z�i���\�������w���N�Q���?�R<,o�����<����-(&y�(��<=Q����7���x��(�B��!�kF^w��r��OO>�5ҥ)D�f�6~��H�m�AKJ�p���'XsC� �2e�z�ն	����D�����~�>6vt����k��W�����x\�[5 ��!�Z�_��������x��,۶�S+�N��b�$Y�*�n�(;P�x	�G�����\��R\Nwx��?޵������2�
 ����E��4Ƒ��cnR^���nl�\$oi�ؑC�#?`�{ẍ��l���}�։��\�(T�El2>>~5�r)��ϞI%6����ޕ�/����W�iL���̾��:��j����0�[��Z��uJ��UK�*�Ġ%T��'%O�u;jD��"R|v�d�>�p^�(�Ë�4Ew['�oW�#P�_����ѝ�7J�������op( g}����(O�n#�$M�t�jai#~�A۟�Ltn�S��F�@��"��%uX��
�"��f�J�0��~}i�����ѓ�n`Cπ� ��G�7�L�*G׿7���Kؽ�}JF�:0n. >!^l��
���2?�GZ����c�j�E�>���d���ib�8VI�1��u`4��5)��D�k����5���a���Hf=e?z)��d�
�n!�au�0��W����и�5߸�5�ָO�M�>l�wU /�9�h���YV� _��fMz����E�1�<*t�q��{	ڶG~uu�B2fZ�K"肗��ɩߐ�B���@�M�"�j�qi)a��
��,����2�� �~��3z�'1Y(��@�)+��??�� ��6P�I������ʝݱ�X	��h�����	��U޿1��H��C���b��L�M@�y!� �z�N��b����Pƻ��4��heGo+�m��N�� 'Е6}���K�8,�=w����xZ!������2/��O�R)	,����I6�d*��h; 6!dk�S崽��"v�������v�Ԑ�w�%��lW�t0��NT�rG�6��k��;� ��Ӭ0�6���I.s^&���	IԗxXj99��-r���1���oqڼ�z&����5�=J�Y�[�z��L̴�[�Tԝ�8�Q��f�:e���a摲�j�#/�K��P&6\�%�#�.ӻ��<��+=N;<�Wz��|=a�x6���^�����0o�n9E:�XRVLd�����^ƼYfK�l�v�9/��u�Q��mg���bx�_� �5U����ջu���v�����A���������p�)��w^�)���C#�O4���BV�]�<�x�5�1zz#/�'�Z����)�d�~�b�ƛB��v(li�|V����+ȍ`�]��U��q���D}s�����%R�6��$������`T� NP/����J�,A�� ��7B�z��St)��חs�W��������0G�����^p�p^r�Ԫ3A֠e��9��p��:��ա��y�mX�]T&Ysm�?X��D��wu�{t2�)��x�+O�ۓ\e̦��̋�o���w�_<�*B߳e��?H�����R�V%����+��!e�u�L���z�X�'���ŋ9o��渇
Za29���n�*A����z�F��%�~�M��1�י��.̐{�xaA�a;�;��,�����ѣ��[��7F��ʊ5j���Y��B��}t���	�e�h��N�eex��q�E���/=��#�;|0�u+���4l�{:࣎�>?����aZ��[�+vD944���V�����
̼ߝ�{�~���O�f3Hh$����jb1X��%�� ����9�
 �ܭ��7�O�U�6��X���-ϗ��yc&����A fo�\�3���˓X��ci<B��ʵ�Ŧ�"��U�l:c�u��@��72���3a#�\0**�#ש��bM>�WՖW��$/Yu)�e�/���S+������3��X�~�Tl }3����q^UI�6�4��呑�y��S��4$O���6p�����;��B�V��1B6$�֍�X�..�9U�-��5��3dn���͢Tcs���g��v�ǥ�7����U����(�'<�>�������� �{]v�=F=��	�*ay��~����@B����eÜx�Y/_���5���8y��A��V���p��Ga
*�l��q0���f�?*��Š�4�ZRR25����z|\�%
�W(C��Bx�G�&o�k-�&7S\�f~��,�"gSӰC5ѕ��;Fy�gQ��h��Lv0���g���&��\���ֲ�Hp��
]�]i����ĔD3�-lMC���F��)S�寯o$+6��EʈxJ	(��|��Bb%?��hqY�G<MZ�>Ϋ���܃��ki.��`aa�9EAQR�d\�|Yhl�D���D
ʖ64K�3o�E���U�LL*�EZ�a)U�����<]}g�v
>���~��A�ձgI ���~�(%�	��*Łh�1��������Cj��"��$r_!�+���1�e�b�o�2������a~�2�h@��ge���ڗ�6./t�\%��9�8����Ak��49zu�x��U5G9��1���9Y�� ŕ�^
��F*M0��8B~�1'�x�"�/ީ�O?B=ϸ2�����󖏗�%uAE/Hl��K2j�,JhX��i�����٪� �Ix��C�ۢ����D���y�f���H0�tӔ�T���Y�fI|��)�'i vG�G_�)�c	����2`�O��Y%��L=�={Ǳ�������i[I�e�Sb�e�z��企y�+;�m�d*�Mn��jYW���Od�����:�a�rV�7�[VN�z(��6�h�g�~�<Z$9����e(iLU`�����N7jXjFF�����6���^)G��0�;k�[�ٝ4X�x����B+����U��`Nu��z��c��	l�-�^�bwPӬ���~c�����<_BR��\u�0�cUDHذRuщ=[�d�O�V[ҭ�����"���Wv� F��Z����Gú��[�{����,���\P�AB/����	�K���!g!��������
���/����/��3#8O��CPJ���w�Ѧ����~H#	n�NOt�M��F�n��'"�^��)��mn���o��y�6��%:=هm�+��<	���_z�!ɀ��N����Z[:��c˄�.i
����7�%��Q�U$��e��b~yg�(&��>̔[2+�3P]����6�n��bR���E�������o��0�O�QYۣ�d}������+.�O~��N�,	��>�\to;wA�@�HZ�au#Q�9�(.[����)�7������?䃤r���<�S�R)k�J�AO��/��)R�ڑ����D��{dϣ�f���F�	3��|<��p=�PdC�-�$�Se�*w�= _����x!G=)�4�0N.,���D;�v����$H������>�p�KP��>P�#��r^���*�,�#�t�-f�-S b��ҁ���l�.c@¨��)�D�RP���`<d!���?U6/x3��[zZ�~�n�o�O��ދ�O�$��[`��*�R�\���\�Vx�=[B���`�f�;���FǦ0˿�e�O���V����Oxl�X��3�504���W�/oE#`_�\ۂ�{�J��T�J�O�I{�H�,��P�^BK}���䴯^��,�~KL$��vN�H���@�z�&�o?v֡���?���p�"����k��
�`� �T��l��4t)++�>ΐ��h�b~鲪"�5J��h?���4-�9��F����莃�#Ŵ�	QHB�wQ��qNb����[?�D$���wuq}s#�琰NL�3�=GC!'ct%��^��2���h/(����	������@����JSud���$��	�eavJQ������};o��W�c�W���~�v�q�_�IGp~�%$�9
?{���Z%t��z��<~�j0��X�/C�`
��R������	;�-�4*f����Ɛ_�Љ�����dq)%!�~���߿6��ک��u~�މ;6ܟ[�l�_�5��m���W��9B���Z�@}��q�����b]��/��9�G��V06��Y#>.]#wrG�*���ݜ#w\�9ee��C�zqLAV$��;{ĸV��IM�u0���M���O�������?:	�hH����JΓ}׍�;�c�AjM%�%h�[� ��9�|Bg�9�[���+� ~7�64�"!o�<H�	�a��.۝��߳UL&v��������+o��X�3tTzA=5N�ʩ�������S����n.��7��'��n������dm�L����cڴ�)���<�����Cy�
�h��� T��}&
��ccc3��8�
eY
��Kx��>���b�_ho��{�$��Ɵ&I�_p:�W����B:?z�Q�� �pE����i� �S�\�T��B�Zs�P��<Ë}��+���H"OO!�#eK���7S�_2�r�����t@@`��F���`��V�S�E�9y���1�������华G��^��O['4�e��S9*T<<�>{;fz�zi��r����$�as��[���(����&�n�d�V�@~����q�����9���GV--Xo}����}k	��b��'7σH6�o���c�Ȁd�:0/C�г72[��_:_n.G������*�������u�Z�4�9t���g~|~s+��rN4~<��P���N���C#*=�/M"�����3	�����@�M����y`��=���T�W��>���9��D�7�-�0O��RM�w��������NY^��2�ܓ)�u{�������{�$[���h�{�=y���핯��rRldLL�@"����y�+0.��>�� HQ���}2��x���!�͹��G�P�ɥ*� +�K��6�B{�	�ZZZ~V$�ġk�EFb���*�o��[��@gda���?�񑑘Rh�:��{S+:R�үx�` ���BT�?�@��������o�j��OQNO&���ԋ��(�-�'W�q4G����^����[�yR�U��i�v�[��
�2�c�p��[�6��dNpH�/��I�rTr�noc�ՖJȘ�����;L�B�h�m�߾I�۳wU�� �k7��F~Z�'|5]���e=^}����? ��3��)Pݴ��I�� ��ݱ(�b�;�ҙ�I��ġSӂ�;5Է��{Bk�Y_}��A^w-��m�t����V閆�/���lTYO��[�<���?���z�@�ڬO�C�>��c���Ѱf�����`�p�"�ɪ���l��,:���*8uc7:�(`���G2���6L�&}u�ż�&JVz�5-��.k���#��7��.�K��{�$��Leahew5����ϔ他�;/���n},�PJ��/�m�.�e�q��y|���wfD���X�
��Ϋ��ę@-�b����Þ��%u����%�sD�,(�m[�/*�`x�75�{��\�p�@_�F�X�H�<Ā��S�	/���i�Z��RAx�,�k���j����%�QK�%�>w��z�E���H�����ӆ�E��E���K�5X ���H:���z-�t�[ްӺ�jC�[׽�QQ�P�%Qt� �3����߈��o��%/���7_؏�+'��tӵ�{���*���,g)<}��eVc
0�(��O��Sl|�|�|�_�3��,?�E#�Z��؃��/���_�	$��F���~��@Ң������IB��=XH����K���_֝�]t3+
�Z��g��Y�Es��;�Ԡ@�8�m�(��tF/t�R)�FU~�;�x+jkV��w� ��ksp.5���\\ja[EZ��:JkRxd'��p��k�6�&���-�H?QeM��F�i�R0�H���<���4�5x�ɽ�o)��:�8+���(�C�20y�a<a����:B��ĥ�"pK��+BSQ�R|ʞ���� *�lj�6��-%�Ά��ZZ�{��/:�����\��NU\����t�.h��r�H?�gj͍��]F\�"�U][r_X{A������GO��ڝޣ��B�*,/�Ώ�N9���[-�MK�n� W�
�iq��Ϳ$m���V�Ƚ�{�q�c����Vc��h�uZ,?��y�doY��c��/�fI�k�5����188�\���2'����Æ���x�6��f��߈��p��r�*/�]	�,�B���/�;U0Y�腐s]3���Pdg	�_�����O_�sS ���L�|���j)߮75�q��8��</R-�9;e��Ͱ����β}�t���E�#�]��N9x��MJ�e�t���օ���[NQ(d�a��ƠH��<�>o�!�p*�'\F_r��P
W��l%w1����M�d�'(K^`x�B	=�b��$�b9gE&���^tsv����cU��2����G�T��a��'̷�;�[�;B�wr����q:F6���!mK�R�+��z,|���C��{r���i���'M��z�
^D���������TE���gY]��2>8��\%�_�b�G�H���N�EBA�cf,fD��x�C���8�iR+g���H-�D`"S����BR/�gA<z��"ު�'�H�i���X�3��>�!W���29�� ���=Y�\����1��� �zÒ)P-��������f 6h�vT3�HǤeռ�h�H&C Y���?�Ƭ�[_�WX�K�mD�;{-l3�vm�Z��W`6� spZ�e�
0G�*��ͧ��Y`��Қx)T{`��e�����X7�	t�����X�Ą��!�u�w?����у,��ìs����n.�7��ߔ1�Yd��c$��f���$����ؐ��^��!���m�Q#��Ƈ贔�BN��J㫟b��ŖD�(�Kpⷘ�g�$�	��,Qx�*��_�����'S��نr��C��X���#m׍�<Qٿ_X'��9������6g�v_1St�P����U�/�'B��A��ц�^��2�ɲ��ý̪�t#�h��v�u2؇�o>^���5��NL(��9R�������
j!�^�|;�4YO���D�'�v�P��٨�		��8�֏}?�r)3ku����U�J��hjC��`�0I􎎍���t�ojY��٘>���3)�_��˝�Ls��56Ҭ���y1�o�q����+^�FH5w����������f$����j"��LM�.�ڵ�mo�lZЀ������S*�q�y'�RaOG�S�p%����f��m��t��x�&2�3�vr��E�т�W�c��rVc5�S�C��H'�k�ЖR' ��2b��a���z杭ٙ������5^G΃BB��e͘tƺ������eu=c�l����s+���� �F%%JYh_#=��R�֥wв����r��3�I���`�VKٷ���β��9�/�{ae��9_�n�nK7Zv�
o>�\4�]Q�5m%o�='l������'�j��h��P��д�,�-�^��Cc=Zj�3���4EHزx��-�WOu��q�WP�z��ޑ�7�H�����;M��&�ltD��^Oտ��m��)vj55���a��٦��["�iA��1A`L������+��qy%-������]t�ˢ��,���2��)��L��=`�x�Ԁ�WU��>�P���g���p�^`��.�F����T�YK�{@(�Ub�׼�"'���OJRB]0#6���6����	�IS�ϲ@?�LK��h�r�>�+/������9l�t��D	�V�d�]�eb�#[	B}֋��-��J6��j�\yɚ�M���j������d�Z�7א�ג���Ȼ�~��[�_�h�ww�?ݦ&T�2���j�ăھ5�[6�͌Qx�Y?p:,��7{�z��ZɌ��]Ak�m^����" �2FCY�?�^1ӊp�ǖ(0����1�$r�̧��l��O�|.m�����&��[�Ac'W��e2b����>9��Y� ~����'F�_�1{��7W2%5`k��������7�?�L4�Ns3i�5�q�ޜ����/�@�<���J�Y�D���
z�o���Ϩ��#F�����������'�Z�s��<�?�IP�}�LA|��H�H+�YBa��P.����­��# �BɮuZL�@8˞��\68�x�*�Fw��N@��z����06��l���vR���82`]-!����y��H̪����H����3^D�M0�Y��^�����P3�5�����C�Q����$oP�uU
����avb������b��ٵk������� ������n��2���aWW�ֵYSU	a�z!�)k#�JV!z�-����錗
���}��T�[-+��Y�#)��U@�4ݿ�yC�Ҧ�� �2'���&ZW�[����eI��8�-E���Gf&ۄ;�PC>���������(��*k�#?��aW�\�q.x��x��/8��/�ᔵvO�/��)��w�s�/#�:2�FHÖ�f��Ux�Jա��ōd����@8[����[���)1�1ws�����>�[	��]�E��@�d�AA*L7_��l!i�u�b83nZH$j<�P@��������y�YeS�=z^l:޸\��<����:�-7�WߟiB�����E8���׬�>2:2��r�+<up��9�/ݮ��b���8ж}8p~�ڔ9=�7h�j:��ol�ixX�x����H���7z}� 6r��.6���=p\5,�4gh�,*����������J$d��U���ٞ��LȀ�VJO3��j�Gp[,�a��ݗ#��`�f	�p6:����l�5蛅�,$!-jJ��;M1AG�����J*Z���Qm
3�����4A����k����)���K���#L1!�CZ� ����}A,�[��$�@��~ry~�SZu�~Еr΅�8��Tc��x�͜���%�Xz��&���ܻ|c�)sw�N��<Be55�QV�C����G���v�ӂ26]޺&�.|����91�F~KKs���%���G��Q���ot��c` Gn�E[��86�?��7�^K���54ď3��ւ��_�=�Y�if�Z}����h�zב��'�{�}0p���܋?9�lu�_z�����?}1��Ŏ��$_��Qxx�����$�ZNE�6ǡ3����^�m��ة�[Ub�"�ƶ��$����!�e��]e$����.��������F�u������K�Si�Q�NlY�z���-���	�M� ��:6��6���r��K������փ�=k�/.����}-]��mz-6~���9�~���60���@��<��ˁ�E�ڷ,�#䍏�PCW��⬢mO~�(\-Z�Dƶtez��W�X �=��NeS�-z���Ѧ�:;"]%����]����uIjVa}���V��~����-���˕D��y*�<vW������ZԜ�$���w["~`�;����`rG��q�=H�]��vAmk�[�{q�Jllm��M��6듙;�Ց�dL��Z@���Iz/�0�k�?$�cܬ�a�ȿlE©D;��Eg��%aOĦ���'�J@�#�mXm��O�p&$ֽ,�.�<	� ͵N�?@&峓`͐��c=XDÎF��~�INv������L-1��a���+�&:�oٟ�.�rNg��A�Cnw�$^�Z�pW��[G�hwpқs����vo�+�׆$v��b������l��	mą�z�8��#�WU#iҮ�?̻��f)]K���IKQQ�!�W,���&͢pǩŁS"p��jE3��{���a�'��+���C�ۓiy�F�n�ɢl�AaSTt]Z�>�3L�d���Rt3l����	���3"F�t�g�7a�̲m���b��E����q� �
�"��IQ++ӂ�7\��ܘ����͘ �˃��͇C����D�1�C/x$�=59��[$�̅�E;��z��=��PO�+$�OP@1D9������/�� �1��j	�lU4���l��N
�X�rs<�=��?r}�kh���X���%��$c&6j��;���P=��y+�_�}�'{����[%��4��XJ��f������_k��k�u��%B�o��յ B��>�	,�VV��/r6j��������ӛ��u��j���r�w���mMo��^�/_S��Z'�'�LT�ۛx�eI���ȳ���y��+S:�t{�����{���*6�W�G��&��9�;��	����ϿW��w!��O	�8��1��C�P�|!iM9f�\�)�\{�@�x<�z.&2���ywb�4uAh�=����w�]P������z/ t� �!~�X�����oeŋX��8���X�fw���'�`Ԃ�%��܃n�c���,�vSː/�{{�OX�W_T�D*চ�Zs�*�F�}l:y�h�E.u�M�#~o��@��Ç�{�{���0�kT��Y:�lm�I�F��b9�5@~ϐi���.M�8�?H�1�If5�������~��d\3�C�a�0}x���樄+)t;*!6��+,��������j�%%�����e��l�sNp�0��Ȋ5��=��2�:1XR��׼}B�]>7�K�/��fm��Bfnat�E�g@�Ġ�Mmic#��.�D--r��9׬�2�8�VN2����(H}SS�R�q�G���
�k�ZP�S�i,��mK�y0�y��s���{|A�Cݷ�&C �?co�ѫ�L���=�g����SWa�O'�tӡK�.����0p�[PѴ�����-2����T�C!mAP����G���� ��Bb�U����|ڙ,�|�"���D�_��Z�8��4������7�"*	�h�F�Gjÿ��w|v�Тp�$w�Њ}�đ�==(L�G����l1���dhܚ��+�9s�O�D����|;?��Q���Ȅ�eM����i�{�T�)� R���Y�oe�T�:���0_�K�d�o�KO�ʎK`��Iju�� /�e���V�k�c�����h�_$B�ȏ�/�jJW 6��=^�n"��%�V���'�`��}�l�^���ԋ����%3)���X�&����%���z��J�jI���=T��0F]�l4�߿c�� ��Jj������A��%t�'��а�����iBWWWJ;a�Uz�z�}���+�-�j��ɢ�L)SG����=�|
��_{5��ٙ�f[��t6�2��Cr�����lE���Is��5�q	Z�����M��š߸����\���G�o�>,}#}����gJ;��llrrw!���HΨr�/�ˍ�S��IC���@VV6*���T�35Ix;{��D��|k�3���5%(��Nj���[�X,I] �s�4'[�tT)rii��m�q��w��"
5Z�f4�"
���Za9��f���Iܿ�"��=m��Ht���}���m!-��A��5Y������Y��[0&�>V�� ����y���;�J��=YU��"
ZF�2���j#�bܽ�Sd����.��(�88,<�U��"YR�Z�^��[uu���+�ϯ�F�����H��'@qT�|/��҄ʊD׮�MJ�;�Tc�X�y��1��`�;�.H�:H\z(~�����Fd:I�;���A��eʳcR��!���D����I/�d�'uʳӭ��w�r1�K�k٭�������ַ��Y�fWފ�~�K����i��S�`zr�M[�1����_���3���lՎ�^D�;��ǧ6���~��m`�_�H��\ZE�f�r�,���,aUCèj;��=��9XXXJ���)5u��7y�,JœF�ŏ���T��y����m)��)\�HA���ɷ�002b��:yI�����y��($���R������Af��9�'+9�4�*�~���Z	�k�����f+���d��L��ˆ��/1#��d`6��(�K@؎��Y�(�a�*�r��n��x;"���SmOU���`ϖ�v��mP˗���ouR�hILL�V�5\i3�[0�$�~�T�c_	&[�C(u?�{���/�h��Y@D[��������>���)@²�c�~x���/F��P Ǐg"q'F�^v(��\28���K����Ί�*�q�￹���o�	�

�jkݝ-���>���/���|,nt:�D�N�����b��3�5?F�_)@w�F��[F�������N���_a�����."�g՞��ǥIc��}@������.��'��i�_-���񅤄��Xh��A���Q
��92ڛ�p��d��/�~a�t�a(�^fT�n�O�1�Ϲ`:�e����D>�������O��9�nԢ�}�֢
�����35Й����rH,���^�d�4�|kf��x��_Q�9@0�j��t� ��;�ʪ��M�R��}ll5����dWv-�/S���Y���3da1y����K��o�{}�a�]ͤ7��1������?^F���䄄5�TT�IcS�S�Š����;/k�USS��굤�RcS'�I5q�}����Ì�o�ЁV��m� �~�Nӳ���ǟ�����|�_WW'����-�|���ݦL�����""��Uu�)�7p�.1&٧$���}8Y�<���m��4H�J PH�m�;>���f����[U�cґ޹���:y�׹���6_�ې^_��a�'�'�_�,~zf:VѢ�������70<6��V������_�ȡ=芦�VX��5@.�i���Xr��P����lj�OWO��At�B�����)gc��t���~���%{�"�6G�:�˸���2[֤�c/�/˴G��{����_��_:Y7�~8��Ă�S�"1!w�`�A���U�3��)���M��r1�
��}�ǋ�9+P�꽆�vK�2g^Tﲋ=M�da����}+�5T���Oʚ�Xl�^�*|n��A�&� �֛B�wpݞ����\����UG��x�e#���#�B��̢F�u.Z�����Q���1޽V��Gٷ^���48�P)z2T��t�]���)5�\�qS���/�r����)����v�T_��ٙR����d�p�p�����5c�c�_����|��ꄏ������
� �c@i�=/�1Y#�N
��I3���*�UZ�(����OD�� �^�a�5�ߙ��ـ�r���V�]�j�'�����0�A)���C����V��%����� �����_̽l�QB��Ϣ������#4������mG"�����+�\��m��g��\�^��kݻEY5ȥ�	�1!w��9[N?k�a�=�x��4:o�VE�Ul�{���8;Ռ�Cc�rooW�g#��Z��[5PZ��ɐ>-�>	J��8�꒒�;��|6z���L˓|9rH��'�I�@]u5^rCC97Y�A�*�������VT��l�3��ݛrG3o�;��s�?̈́����N0Քm�6�+X��$i;<����a������4�I3.b�+���xl�	����OF�*�<�h �`.K7mt�o���wz�iI��ʛ+�Ρ���� ����Ig&���P@�Fԯ�ɏ����7eⰰ��t�7ǽ#����,��[[f߮��&�#C�γ��ޒg����x6m���BxO�Sβ�T1P��cߓw��.Y�7nu�)*�"ew�f<@��}�}<œ��|IiS�d�Ө�q{fL�B�ŉ.u�x��R��ג�O��k����/��oP[�D�N+��������M���X4/m�ܙ��v?�'D�Ğ[��Dtε�~�=ԕ�<��iTWd�fl9��#���_1}g���F���&�����ϬQ��_�<`,3a���ߓE���Uӭ�=I�F� ߚ�⼮��5�Q�����"��r�a��ne��8�b��NTM��/�Ċ�C.	iy��?X�qS�.�p�p�K`�����+�(}�9u��R�֑QЇ������/*�]���� ��|�m�ܤt(�\,X�MUmv'�eg��Y��C�#�T�)��G�o-��=iqY�"��������RV֛�l3A[&��3n�KO��S����9l`����Δ0B���\V21��^�B���@ddS��=����
����P\b"	���2�h����|�к�僓L��`3a��xU���c�Ne��X�t��z<Y۴Q���Y(��B�ټ3p�d�q��}�~8�+��FFΟme�|_퐟ȗ?{�A,r⢣�\cC��VF|^�����;���Cֺ�S�wi�亍�q�ڵ��k��ݼ��jM�6Ir up]��,mĵ��S�H�����`x�;�u�Dzj^�����iO_�?����YRNJ¾��6XNᕩ�5/�"o#d�>a`+K�ؼ�Q*�bi�*��.�D��w�Dw�w'����*��P�emEL��[�=tc�ҹ��O��u�ykލx���:����T�4dG�wH#c��Nq:/I�Vl0�����IT?�MvEg��6��*yo���;ވg)%i��~�<8� 
t�:�Cxm�������[7��\L�=��F��?�{u�i���<��c�mR�t;�b������i�ٜz��v}��櫌�I�^U8�eݑ�����aN�j�>%%���a������00sp�m1��W����''k�nC~���F�d��J�j,��,���饧#��n�
�=���1�2�W���O-{����^���"�|�'���6��R��)L4�J�-�����m��v�xx��,&nQ2�T��$q�ru�K}C�P�<����22p�YVT6GM��_9֣�y�9������������_��=���s4^�ϔ�j}���y+#';��V����-ǀ�����	�E��R��f�u}_�|9�B��|������yA��Ϊ=�+�1�T� �ۘ��y�m�JH0��ͮs3�Rtj{�3?�G}<�)�X��ԜC���e�mPW���p������I����#�㠎�?ك �_��WW����ϔP���>0 7�P��1u�����l��p�3�jP�H\�J�$��`�d���PPɨCS8ֺۏ��C��}+�т��j�*��܄I�:ó�ޞ������4f�v'�R"�:�������ҬN<������~�c��ĝg���Y�|���i[���}��ǣ���b�cɝ���y'��gG3-�	3V�)��?:n{��ƒ�eA'S�GY5�f;���f��I3zZe��"����4�)�<�B�����(�0:����FR�?�za����P�T[S3�T��O?L���72����5N�F�Suط7_�Rt��^JJJn�7TAj\"�����]睏:N��/88�Ԛ,�̿m��rެB���`k{�(��q�h <?��U���R������Ǥ���q���	)�+�{��	�.V�Vw��Z�B��Gp�9OV8zHddtfza�&v��)^���G��S9��?c*��N0n6�6u��>�	�>��"���Ue�,����}��A�;&�k$oX8Xb݇U�C�:���3�ƣNsT�>}��`v������Ķ�s���Ox�	�5�˳�u)x}�a0�#TLs�_2hW�d��+@k<b�.�����%����C�c�K�� چYe�'�dėb7�q�%:�(��'� �c�}���7<46�Vろp~��OA�*�����HĬ�0\t��(rç��ag��x��\cc�e5�PIG��:Eȕ���{������«	�V�3C���oqqxw�NL��v?Ĕ�p/�w& �L>.����g�r��O�\@�Pb�JB�+��~�Ĳxr�ZRnF1#�е�1�������bPo�o� a���T��b��j�������z��t��'1�����<Y�����J��%���C��3�i�>gVk맅f�{��Ͷ/�0Q�XU��Y�$����{<��������66�A�}��ظ8xT���c�&W?u���3B ��:5Z�U�$�!6=q���)���#lG�x�S6~�����)�]&u�tX�ԡ���i���x[w�>ܱ��~?�(*���a]\��ϒgg��wi� @�i��[���a�U������$0����5��WlAn/�v���5�H ����;)B����C���Rz�Դ��Xa0����n�����v�s���IGP�0�a��̊�Ѵ���3ס����f�ffE��͗K���KK-�[i�k� 0:�V�0|}6�U��������^�uM���f�Z�	8�3ȯ�C:�����D�1}w���3�&���c!�����#.���6��G_�xߧ�G��Z$#���'Sj|�����0����>)w2u�
��<(v�Ʃ6�zę#߀�r�|�D���=g~�k�#�a��	�����L����Pё�'iJ:��`mz�׏Q/e\�;�N��|듮p?��~(���~��S���.�9����>���)�o�I��G�~)r��`?"<�4k��%���u�m���ظ�p�PC$�L���лݘ=��Z���|w��[Ȣ�A��L������Q��QQ?_��"�% ݍ��H,�! ݡ�4J�.JK,H	HHwJ�4HI7+����.~>���w����ρsv�3wf�ܹ�ug��;�{vJ�v1冼2f���I�Q�xs�&�㷎E�ի�Ό�/I��o�HB�%3{mIVto�|��+�5��'�m��H�KZ���P%ὑ`����G�$H��x���yb[N�l��㑨�w�>��2V��w:gFfv�a5�v�<#a����}&N�p���;8������d,2�̈́|W.���CS�*X�JgIy{n��uf2�J����6��Qx(�.y�̪�-��F�E��{slfo�0S`��������t�[���pL�b�,+²��Cx���M�V"���7�n�����͏�f��Xm��=\�a����zG=��n�h��gA��9�g'uәOq/[�Oz���VB�	}�e��5�X!ll��f�ك��;��x&�}a��,��/d�$ȅ�.����@=�~�<����58-�a�ڿzV@�%�W� o��zo2ے�--�'�����V!�g/�,z�1@�7���b�R �O��s�У��!ߚ	�H�9y���7a�ԣ����S�>�Aב�����E�U��q�"��K��K���ߪU&O�@~#;��e �R�]6ceq��7V,��t��W4U���`��٬���q?oJ��>��?�/Ý[o&�g�cK�:-�)�}u�kι�<���N|���Z"�B�Ta�%��!�z��z$���zp!GB��#�Ǹ�R����Bv�b��j�<���
���0�4�Y�_���[�u��X��8��������l�r_�TZ�J픵��9�NWb������ �Bx\�Om�فW��eKc(@�� [�װ��o�_u�rη��A{���H�()�q+>�6�#������<�I�ŪK\!�y�{H�_9Z#�G�� �G�����DP���-�gZ����DC{�=N��)����!;/og���uSq�Fd)@~��U#p����UO�m�E�iY��~��@{���=�q��ŷ���>��KD;�`��ai_���Q�GD�'�>*�c��G���.�@�9�Ͻ [ �,V�y�� |G��ƇGG�G|��L<�S�?Q	2��-ܳܵ�^w���q�&�5}Qֲ=o�����E�r�9ǡ���+���V�-q��AًV�y��c������#1�)�{ۦ�|!�l�I1#�=�1�U����FH��n<����?��B�1l�#��%���J��$'䊤��~�k�G��������:���n�и���*��2@ ���}nג����:���喫���?�^Jm��b�O�y�Z[W��]"���m3��Q�3!��sA���rX��B�v���������.ȟ����H`�}}|6T���3��r�8�Z t�(��ϟI��$Nث�)���}������not�UA�YOn��cu��ˇ�ק[o~��RU���=�d��������(�E� |.� �FR#��t/;Y����/�J�)bP�WM�GC ��M�����j��q������*<��������4
-:����	U��������ɍ!ɻ�J��`>��L����[���$PߓH����fR^S�G�B!���7�ʳ�e ������2k[h���G`<�wq�f�;C�s�z|�<?�\���������h���~��r�ߙ0F��#y{iQ�e��o��r�)���ÇU�\�
�a��@���w&pAJլ�KO� ��R�n���l+���Y,�.xFPʹ�#�[�4�V?D}Sn�{?ț�@��z<�(<�3�W�a�C/��(����L���򡞬�Ն������o�g`b���,���=w��6y^��s�jn��+)�y�5݂�������N8)c��a|�6r_G�U��{UԇQA���:!���9~яb�H��->��h?OP+4(�M.��qx�>���4I!6.��"|�=����<U�]B`j~�$���Կ�X��ռ	���P:����y8��\��vB]bM��E��w�n���wD��~y(�z�zA̼p�4X���y����	Y!R�O�E1�T����}/�BB��l҅)�#)ќ��c/H?�.�Hp�U�l��DXVI����;I����c���!vޔ�W���7�:��u�)k�ƽ}�Df��	������[m��A3��*��[T���z�~u���nnn�\�����E����=�����%�p閼�f���
�ޏ��-��B�.��LMݛy���D���ɾ��@���D{�m�7G�0��fь�=�-Iet��>��׽�r,X}��\]��������LϦ;&&~�ĳToZ�~��NX_���ү�|��������nY)v��ճ<�h�f.q�E5�d��{��ȉw��燽q���,Bb��?���N�����؏�u�U�ttH���Ǘ��@�p���v�w�n��B����cRSK�}.<\Y�[�=&Ë�5<*�@��B��=nh�X%#��lP{�a4&�8O��DC���x%׾L@���D��VB����ʹ�m�"����#�o>�s����ӄKKK�O��p�śUA��.����OE8���4�w[@���M2_:��I�����_�=�۝o��~���I�:l_i��7�Ó�$�G.uBo�9A�'qB�ޫAM��O��lxJt�W��</V*�W��������ȷ���VV9+K�VV�ET<I2�V���B$�:M"��M���*8884���.:4AY��0ħy�xH9�����ͫ;��FE�PM�G�޲���؅�����]"u�������w\�c����f�qa�c��6+[a3���ȌD����VwdN����v�*v7(�<�ړ����NF��SL-:�Gz�4�=i~ݙ�����&�o���W�'�g�=V�z5��|�L�'wF*Ґ�qխ~QIn�X��x�bz,���\os�6Bk,z�^�>�񃝻���k���+Uێ�{��sKG�J	����I�C���22;A@���GMa�8�3��nB_ƾ��1���M���=o�&p�Dd10/Wܰ�$�X�"$��%Xj���y3�T��ؿ6gzܸ�Dqy���>�g�AR$M7��95r��'2<g�ď����h�
]��8b6M�KP��|'j٧��(9��YZM�͔���d>�_SO��E;LI!�u��̾I���²9�i��H��~u�Z�sY9��N��1�*Ff?U�8�v0�&�;�����v��Y#������>��Ä!���?�;�Fڝ��͚U�����(i�|p�Y��"�*�G`�R<{]���lr!��Y�'LV?m�C��������}N.aWK3��,�v�b޸5��a��TT~\w�3���>�ˣ�������ˀ�/>.S����^=�ٹym��zsuև���6��g�S����3+rY^�0�Pc��͠}�z\y����u������vi��ا]YIC^�A�S*���ġ��3��4q
�w�o�3�v�S�����Ώ����Y��Q�G���]���$o(������	^�p��P������<����һ�B���#wro��ͷ���xw���mD�0���0�������yԝ{������$�h�ħ��ta
&�y��[�R��)~#�1�vԆ�}c�o���J2:K���L�{��2���7BMS���BY�t��7;�<�cK������r�ϑ�9����Z?5�m���	@�k�f�)���NH�8]�")9x�C?���a��..m�[c/�l���=�V��l�r`vT�b�O6��Ӈ���%�⠔N+��=:�3�|�?��&b�#k*�S @x}'�f����u79�0J&o���1�����i2�֘*}��ڦ� YZ��m�)�\�s-�� � �3.��'��DF�
Vw��%�;�.�B
VLv�~�.4N�L�P.A<�><	Ƨ�hM�B�I>�Uŀ#i�����F|�������b";�ş �I{2h��C�⦦LӔ����:kS��;�?�M�
�]��(;0�0��ݞ���9/�)�P೰���G9���J]]�3ĉ��z�pEso�fH�r3~�ψ*��D�\�N.x@#k� *�xe(k{µXB�k��4�H'��D��5��ہ|���w�7k��%/N�$	;&��ګ�/�|궭�e�4��7���9YBe
�q�_5�a[��X��3���]�:Ch%��o4+y������gOekު/k�J$`ѓ�K�Z�;i�G�/VR����12��f��	�'7ޔ}+ܶ��\N/���-���/(@����w�t�-�����LT�X��HG��0��W��}�~Aee�"�		�;77�|[|cy�g�G2,~��]&d��+K>��z�4��Wr��ؖo�.�ip�� ;���c���1�'\
v[�~#�y���d���Mq�,�򊻛�~�?��˫��\\/[�%$h�D�:���#�C�*,�TEq���k�Z.H�?4������P�����Ȃ.-j�P(���h�7����А�⁷l"@��R@?�Jg�qQz���K8t~f���U,L�^'^E3K5������҂m}8G�L�^�y�^�
{��z}ڕ}4E�C5] G�m\=c%I7O\A�����G���O�EzT?�qȱ���-9F������et����Ϛ��.jɂX���e�M��h{���%#m�JS�u5���h,V9g��4�/$M~�#�Ɲ��������mM�1ͫ%�.˧O��pw�i^q;N� w��=�ֿݻ#��v�:��W�̟��&�)+���zc���#���#���o9ZS�a瓩 !?Y��H�@��I��ljxפ�}�'1&�ul	?� \�=2�qH�P�@ծuH-�=`���rn���A��������|�i��9�(9�G�0�&n�Y`�����>�G͔hY{%?�=ﺔĀж�u2=+�5\��$L�F��e$��\���ϐ�f7�����%�h��/3FW�3"{���)�A��C�����~���^j_�d9�73 ,�����A�t></#�g�
�~�y��x�[���d���z��/D�Q;���#Y
+Ad�?���4m?��8.���ɼ��e�JGx �X4�Y�7r׸��}���'�6�]�����^pF��t@ ��>\(}@�vC���N �]"0�s�w�/yE�d��J~sq�L��mY
1嶨	l�|���@w.���I�et���קse���Q�yۓo� @9uTh��������ʃ>NJE~9>�JD-�sZ�����˗/�GN�_�uuua�����>ddb��M�%N_k(���`J���
?gP��;�"��̂������Z^Y[Y��|%�)P���3v	���~��E@�ʸ�*�Q��(�F�a"nS�a�cgI�Mvr��p�ݛ��@/.N}�gsk�J.PU3��?���뽅��X#Bi�ˣ�ѧH$>��)��6��4-6N����� �\9o�>/[����0Y x�{ڨg�UV���1�CGu��T�c��.*t�3�$ߍPLOI9�1r��fjV����RX���
W��z8$�I+�^,�7�MEå����ĉ�y�7�3H=�ۦ?C"�,��V	B�"x����W��J�u:�Ce��<Whh_[W��~FE-A�����(�/��-��翏���T���43��,��Ƿ7�6އZd^?���n\`�OLUW���ur*�lp�+�e/(�_�!��S����;yj}SSK�;H�aV귂PFL�-�	��vJ����w�tE8j��3�\5���Z���G��������K����݈�H���'�X��	������eY�(M�����C��%�AK�s�����%Dp�M��[���(��=9�.*�벂���dy�Ŝ�}X��[�|�d	2�aRT�"u������t�
�"έ;��b��l�T�ck�.��5_��f��]��ax��/�������`��׃�/���G�P�+�x����dz#�6q+���L��W��k�q�lv(�n�cs���֬ͥL7�w��vx=7�gW/9�'H1A������e�䚔Y�d.A��?���s�bBg,�j������΄-8�~eۘ���6x���,�O6%s}�[�6���=svI]D �ú�0-������x+���5��d�3��%�HJJ^_1�f�H>���B��Uu��7M������N�����Fٔ����m�H)��@�'*�)h����B%<~o��æ���}@�l���|�h�(Y?�{��^ν켖���x��J�bK�v���h�̩��m@�	�|�U2�w�|�M&��6.�B���$5���s_��e���0�[���%J���&*Đl��������/��&���`2O��E>ͫB�W$!�a����<&~eZ�Ҝ��٩��ď~�6T�3Q^�~����L�Rֱ�S�U�1��Hdr�8b�%�Z)���,��lF\<��~��x˪?^_�y^�>�RC�/.>�6�S�s?ළ=��9���>��X{e|�
}�`j�H����{0�����>�e�a���[k37�+FF~��.|�ْ�@���b5�E��]��:������d)n&1^���V}�I��Xy�L�7+�x��?��%�%�i�C ��N�s
pÊ�z�·uw
��8�EZ�s<��լ	��"y��+���S�{��p�=���{:���_n�F^i5��7�}��8�^��e���L�����lU�I�[�����mƼ�25��)M���4RQ��F�'����e����݀��5�+��أR4��4�s�ۤZ]��-[[L<���z?Hd�'~Ә��+����^�<0�4'��+����q4�0��C �~+���E��:���􀇎Ⱦ<����|Q�m��u�8�GD!ṕ<�}*/6v�mt��4a�uY�1�Oa��*N��^༫X��e�9X�{\�������G@���Bk�*���j���r!����yxT���nnG��M�������~�U���:EnZ7�=sc8�gK�h���Mw�4�#k����'眦Fd���ޱ��0������\�h��r�l�m�J�:�\��˘��VH�U�Aj��d�X����v;����2i�����}ӳp<�TZJ>[ܞu5Oo)�:�Ml�+�o��d�|���nW|87gٸ;�d��z��*�Ѯ��Ŗ4���WF|�I�?�7�_�\�&n����۪u�0�*���$��I�{�
'��/����t�by�6�A'���|�V-�WN�---����"���6mn􇪛O�'&��s\��5�pI]�6��4�z���l��N}�3KmS����j�A��:�g�2HL��*��?H�/O�l8�����0uϦ�)�1'�������:���<��qp�=����G5W˚��v�y����pܦ�"����,򯭥�{{E��<g��lye䇴�����h�&Ă'�O��8������v�Q�Y�ojn��e��V-o���i\��ؤ��=�z��^�4�X7`|���8�|K�~ћ��Wp�������y���y���֓f"-Y�:��$Hu���w�Z�����Bi|���mٜFVU�W�:~�Z�î̋��|�_�n���j��~�\{�M�]�:zƄ��R�u��==�Q�r�������r�_`���J�qB����5Y�񮳀Y\��1�:x����M-�BM>3s�6���S�np���^Ҩ����6�9j
�V8\�]Z�q���7�O�\m���/A"�\/~�N�2�9����(q�]4Mۜj,�����<V�O�	U�`��K� ���Ȯb���}X�~��hCsx�O��}ܙ����􌮺_H7'�����hm.4�T��k�^!ˑ[����KGQEE������1	��^�ӃE���Y��b`�g�h�P����K�7��I�S!�Z��#�!n�Guj���IO��L���,f��(�����ԄF�,o|.)!@�4c�,�˧�!Q�b̌`S��g�@�n���!n#J��@7mm]!OZ�5�޾ޟaL
t���2F������V�W��1�Q���Q������H<Z���On��jɝ�]�e���ֱ��V����� �~3QT��i�vzA�g���!"�F"�]T��j���gcz@��:T�֌�_Fs�#|��82N Z|�Or����ga6V�bqA��u����	�a5�}@�[�����ç�����U�x�vS�$Υ;<��Eg���D��rr�����s��_��,mɡ��v���صu���?�٧�_Xs�S����R�����P�3������1����Y�[���@-l��P^q�x��ۉZL����٠��xF�I&�������G��iD֣cG��j_~/����MN�Ǡsq[����0��)=;�Y[�0�dL�1s����L��y��sUn�e��~�\�~-�!뷽Z2؟�+l��ï"�ɒ��ì���d�����	gD4Җz+,�����g�6?#��E�c!�S�b��.�a,����-<�������,���w�{_�.��9�"єۧt�<5�K�����!Z)YK��;��/��k����v�͈\
D�d-����`��[<�O�Í��f�C�\Hg�D��8����4_�}�Ҫ�,�1E���<jFd�{;�o��㮊������cc���8���n�wm����҄�ׇ2QC�} Ň��T�������9��PG'����@���E^�������� !�0�|��D��y�?A���D9ѥdǉ��
�%�Y��ū���3&I  G�ǣ1w�b���szˀ,���׿�}*k�9��I\&k(F���PA1Z|��]���!Cm���N��--2�h��ϟG�Lx������d�?���_و����]cZ��?��c�a|���GG���% ]R�p����ϛ�!o���*����~��Tw"�IS��0��h����p)���v�[/��r����C:�1��C���t��7���O�XXp�Q+�~T�dw�p}aZ��>��7�ޒM�O�k�NN���n��En�H�p���sr��})t|�Ǹ��k
U�&���ѝ��_��u<��߫��є>`S���Q���E�\���m�����^�=�PΟN�-�`VA��F�=�Z����B�SWo��'T7����ʭ��|Z��g���у1�����>C� o��㕁�Z�Ӻ���¢
��Y�6r!��6��*���3�?�ϼ���+��-mni]{���,�B�T���֯85����]��v6u.FO;?��z�����T�X��-tK�p��N���Sm[is��L�����E^)/�}�Ze�I�w�F�N!�,���0��ʳ���r�ׇ'���k)<*���H���T���\�`6:н���CD/��K�5�Nw&�Vz"�l�~�Q	L;K"o5in��1�rAu߃Z#�^҇ms}��(Xf4i�q��w�i��*r��M���������f ��W���𙍿G�� ��;��"���/g������^�I��6�4�!R�Z�H$]W�����9:���
�G*ii�fr܊HՊH�����f烢�A
��b2�`�0���D|��C�����)�T' �<�Z(J��}�݈?�M҄_ͨ����\W?/{�1��+��v����m��η`a����uј���:���辧�ʪV��{22�f�*����G ��
J�%*�=N"OL�Q�`t�o�,eo�k��8�_!tN<vK���/f��K�j��K�"
f-�>]b��d�����nȕ�-1�AhT��73�*_������)PS\���JDZ�s��쾣8z��a���(h*}��m��ow���X�5�%F,C������#���b��ɟT��}��"�����=f��ғ�S>'y�wD��̕�'!�˟�
���nڻɾ+��W�^F�^o��;��R�Z۾7F~~�P�#D�|��
pdӢ+Y�[�^=�
B��䔻�ӑ8>'!c�_����/4���64&n�d��҈�Mx�O���F�<�˖�J-�M���9-��C(��N�5^�JYy<:'Zž��D&1㷠c�v+jߟ�}���n�=0$5��lu�ܵ�����W���,��F��I����C��~�&*�����#��0zϒ�̚��+����{���"u3
!_٢���/î�����oT�S����$��ky�FK�*��ה�]bNt;0�2i$����� �M���e9�L�֣Bc��wkk�Y�$���(���	�h����|U����֓T�<����m�7C=+�G�m��ǩ?K�6���;�So�d�Śr���11>}/0p���X����i������й'z�)�L�]�ٗWa'�D/�)/�_	�-�׀�eKbi�м��֗�t�O�w��~WA��#�{�-����m�0��=�^�Ec�ɸ���j85�]˟ӈ^YC%�{뎬�F��DG����?�;;�p|����A-(��x.��q��R����b���*P�J�|R
�-�#�)ؼ�+�_|���beV����{�uH��*����t{_(�m��-�$rj���%�B�^"9{	���qZ����BC9
oo��E�	�h�ލ��.���#��jﯧ�3UWF���6���ς�[����'"3\��e��?��j�=7�T�q�>�6�4��k'r8)��O�J�.{�����㤿bw���K�L��뭂 �'[M�vq�n����?~�]Ѣ!�\���Lǝ
�N?�{�g��^;O=<��y���E����	��Q���l�Z����E��~�;-3��*G7Q���Gv���֘��V�UI�x��{����|�4�o_�q��`u,g�L��_7#�>��I�B&��t�r�����k�`:U����k�"g+�M}��G ܮ��/��� ���&���+�Bk�!� ��M�S�r�qs����A4�����c}wǕ�oW'F��(�m�,��[Iu��<+8�s�wE��։�H�hr�rݾ	�b��x�ڮ��u0pf�`@���X���,J��u�c���[us��k��¢B˟??��]��q��Y�pS�x0�s�xp��ST���دD9VV�"�s않aO:�Bcy���B7޺m����\�DkRU�|d�:�C���j�
1��U�"A+7HVI� '�Ή���^����F���z�S�)���^�K�F�v��z5�5�9�á1���O�yE�k%�uܪ}��F>+�)U��9]�q��etO_��n��K�t��߂��� �ur�`����J�yD:�{f��ph����՝3��rယ�����U3�2w�B����~��c쾞��H��XGHU!�=^�1<)^���u�Nj6��ؾ�L���T1�7�ֆo�h2���j���i߿�֤
��q�?����q�[خ�[�>1�A�.�յ>��0�Td��*��Ƽo�}����tg���-�����
��|U�S��I��Jf����uZY|�,g�k�-r��*�;�)�>�x!���k�&Zm����w��y���-D0�c F!��]�IʭH9t���'Yh���TQ�=��/b�ߊO?��2�&C�Ё��'��R�,#�Q���Z<���Ԏ�� G����l%	ܝ�'f��L��~��=���M|����7Q�4wʿ`�r��}����T��D��9����d�gZ�=5LM��N���:�	a�\���B+Z91LEIe�W�+f�8us��>�
��G�?ͤ�G�ON~�z^� �Z��
9>��t��-T�zJ�G��,o�"��~>�>~�����Q3��]6�4_$�,Fh!�EŻ-�0�,"�Npl�yB#��XO$uS�(��Z+ͧ-�, 5��ZP�Z���F��������}��mFP��E�UI��\��K_��e�{-^.�jR�[}mOQu rKZ��i��O��!������u�@�"�yHi��f�45q��'=���4g����T���;���Z'k�j���C�gCyR<S�F�2s7E;F��b�4l.�$g/��J�����K�2܆5�,�$X�B�skh�
<��LT�C��,Z��%@䤁���?VH�!>�䮴�'��O���~��[�C��x��.M$�Gf��Y����Cެ�8�"[[�;w
��,�
�L��H&��ڮ��M�yJNB�/����74MC5/� ߛA��qɒ!��3���"b$�J�lWF);wZLk�K�a⩱��]�_�!pt��>)�9�c�ީ�9�@�"-S�&�P"�`��`m�{Bٟ�g�O]��s1����V���x�F��U�
x�j�Q�u��1�H�5��8����c�g����7��P��-n����N��ɷ�W��z�i�-P�A��r�����[}���(u�"{��������37��͏,^�qG���Y���p%x,n�9yk�e���u�v�j~�5�T�_����94$k�/곥U����<�u�������N�����[55t�RFG�r';_Ur�ҐLL � ���D���V�cP�����i����'�ۑT��w��*�����x�W�^ԕ6�R�Q[0[�� ��_�	��y�T�����Ĉ%�t�tܕ{�0:#��J�p
[[�:�t~�Ix���$��J�aR By����LJ����5��C���������&{8pG���bW�	���i�B�/]�lG!�M�R�5����t�N�|�����>�vH��<st��ZO���( ���ޯ��p4č(鿁K��w⒘��r��Z�A�O�
J����I�9.�(EӋR,�X2�Ѝ��X�C�þ� )VL�ە��,ϝ�{�f�4�����g8�U/e�d#;�=[�H9�Yx� ��g_l����K�R�
'��>�Z� ����&�����HN�s����Nu���ss�<ݜ4�iV|�@���`���)�s�32o�b�y��l���%g�
t�9�<����2f�N�4pPTX���&�ْ2Z�V)t��#���/�2��o�F5Q��c�����^�V���4�ل<E*�0c�H�RC��㾣��	єÚw̌nxx��ۉ�y� L���& N�jF�N.����u���s�l�Q��391����RZ������G�l��E������p��v���6��u(��,�9\�4(ҫgJ~v2� 増/��ۗ�,���JKH����"Aro�>6312�\�>�%�#u4���dJ�ļ�5}cc.&����h%�L�k�}5�LpK��#�d(��#���.����	�~��㡼*�0,=$&���O���L(#�3��)��X��+�3e
��y����M���/��>6�#fL'Bo�3����C�95�
3�_�ѶC��8�Y!�r<@�F����%�L	4@��S�8�"]%-�ؿ�7��=���X�x�	���t]퍩|���O1�W�y��	�=�Р��B33ǂ�]�7_�BO|�����6#�.�k�ރGUϥp,�#b�0p ��TTk��[�n>���K�}˅)�&�n����?Z9���=uj�����J�C�4���9��M� �5c1l`V�H���������[��,`8�v|��a`
��E��'2�X��V����U�_������g~�.�j��4��;ri��-Z�J�V�h�͢l���T��'���_�CV76���5�3��/��o����Q�4G�6h��¯։Sd�����|�����B'����bE`K-�{��=�'=^&�7���5����
M���������K~�M�W�/SZ43+�'���RY6j.G��vل�Y��韛����Q�� ��t��w[l�fc��-���>������J0%���w���"BB� @²�~bћ8-�G��MFw�R5����"u~o����D��"��H�^;gS�f*l��-������ј��
�F��(�8��%�B��v�F%XG�iJ���[\���a)��|��I��LF7���~=]=A�J=g0:�{?=D�b5��+����� =�}|�2�b�ȿ�Iw�Q���5��THe��AB�Wjz��V7�~]��Tm9"�V�R�V�H	�����������&[�-\�՝�N1�:�[Ё�:�Ll�E��0"�J�KI�2a�� �{d�"-T}ܬ��Yjb�]�����*�nU��a���b~8��43�qiq��E���3vI�6��Є�,��s���gQ�(�ܭ������">ZI"`� ���NI�7���m���+����}ހ�X���@i��,E�H�����twlHRt�t$��q�6z�T��~	C���-k^ː��1'StS��4�$������롦�L�D�,�nv�t|��[@��-��IB����J�/���R����'At�%e��O�E��w�j�U���������9�0xk4�&�E�(V=�����.�Ci�}���4�����ǹ���%M�S�aKsk�*�إ�b-H�,�����[�݇�`9��ֵ��W�-�C�� ��ֵ-Vח��A�s/�浬��x�u�J�t;�������}����nH���kݞ�#+m����<����
޾��u����W�-|���X6�2rzj)	�E�b�l%�>#m����$�r@)�2#nu~�ծna[_\Z���G������������f#~P�_O+�ݫ>D���|5>9��u$�(.�P7����ۗ]
�7&�?)bOT��f��g��~\���6���.�HN�Z�͢�?��0�r���B��9�Z��sv�+���e���6��D��^�E��+s5١4�9��
����s%�(q�G));{��H��C7��B���N|�٤Q��sx~O\��/l�֏��å�3Z_R�٨�����3�}i3����H��@v���ѻ� ��R^��)���FI񓀱�C+dZ�����|�{����{��I9�\�Ёl����?0�������%C��~������?�n���T��c����},���eͦ�w+t��푪D�.�[X��o�����Е+�c�2�4�Im��E�Д1�a��ݸL�F��c�E���Y���e�����0�j\`r����\k|��J��nL�
	��d�%'):�w}�?��X2lq1�{w��9�@������|��R_X�G�H̫YF��r���Ef6/N'��T}a�Uf�LƖJ�H9�3rJ}�(�����M��F"���7��������2>S�&�����m���ѻ��5�$�.a�RRQ�$�e�I���v,��x=S�[.���@f���HJ��w��Eִ��NM;������rd&�N4���luf~4G��|9Z-��"��؇Ѕ�=���f��2&G��T���7w]p�R:Xln�!�%�:j��K¾�5�xxm�b��\,�� �|�<]�D7zg�={��c��)�D��r6M�?u+Q=�I� ,�uR��^d���<�l����,�t�௽#�!@K�sƾ�9��Kߩ��'����1��Ew�ٔ������A"t̋����� UWS����>k��C�!x���&t��@�թo.+zh: ���Ol21��L'�%.�hy�7��8h����n_&;�M�w�MK�#����ENvm�ħ�o����N�xABR?T^��=̰y��)W��N]�(��$�-	(8�Q{�'�}j�?�<�H��U��np�atj�>c�~a'n|Wu���B�]02{����.�p;c˖fy;E��N��r��yx2�����0�]D��+Ei��%�ξ��
ތ)�Ȱ,�b�zf��2�T��Co�#G��ngX���T AD�-�;B���fm=f$�ۡ�ۘH}�l�Ŭ����p�	��*<�m��K��LI�,�����.d��5���-�єЏ����6 A^��ro?��.��ì+@�!�ry�K�/Q��P��\0�
�̎"���^�/V�*8̪�Ԉ�td�֠F�=�|�t-{�M�"�f�t�(�a-��7!�"+A�����������k��'��uH|����g?�c�zxL���<��E�ѯ|n�rd�W�2cy#�O&C��~|�@���(�_���m��{����&�q����7!�U����A@���H%�??09��+�%��)O�^w���f���������~dަ��y��!"�C�	A�$��?�x����!�~�H2�I~	"i����&7�l5��b"��]&l	
dr*g��;��)(�c�YI(��wO�=^.z�I��,)�F�ѲR�0̡�Ff �ڙ�&Rgp��K �
�#����&���M���ag��bi��@���� ���:s?���R�rdW�=�n�4V�o�m��Q�P5:Y��u�D���\T�쑶b�� �'ui쑩y�̻��q^��ۨaЋu@���^����\�xx̜�t��QrT�����?����X��{F��:}#b@JL~�ЀED/)��&{���Jo�a֞دf�����)��g��$���d�KC���YqT���0���!�R��A���.��U�����?�Ѹ�kU�<�Q�,0�)Jq_��^Y���V-/G�͢}�E$
 �9��p��!�a���7$��Q6����sU���z��]�5�֐p�N��rct��%W�/G�y����d�\��j��#�"�%�y�C�7M7�"�_/�m~��.��M-�0���w]$z}��4n(��C�C4��>���<���=B�8BM�:��fZot�-#j:H��X�2%���=O���7!�m�mG�\*�F�����?�,˂"�uG������N#ʫ#���}���Ѻ;�Pp� �;���9�5�5/8V�����z�?|�y<���?~#	Ee_G	ٳg�B��	�B�}�%YF�,Q֐}���!��:3���{�^�����=��s�s_�9�:�<���gDϋ�AaV?��0��oS�\�vϚ�L$!�O`
��Ƒ�`
�]�畾����9�t�������p��y�uð^-��|,��8nY��-��Ag�Q��S��o&��g?g�O]��	�-n��㴫|�7&��D����.N�u;�N��"����n�J�T-�Ν>\�򲞜#'�4�u*�{R0���,����pfv�#���W0����T��m�D�8��o5���������楝��5l03�EslRҩSOi�5���s��Na��TTuc�GΌr�����i���s�s0n�z6}Z=�8��훬pma�z|k�7�lim^���(��X��H�Ax:�|�Z˼O���b��)x�����&?x�+	E�5{\�	p�o=©�!;��5�.A;i�:������.��̗�|�\�c9��p�`m�[�%�G�Ys�t�*lhy-������c���	��.@*��-�:����j\I��_�ǯ¾��y����Q>��4A�|����� �Ξ�v1�Սa�n6��m���]��ۯB�񵥟b�@�A�6:]>\^�;ș,��j�c���D'z�^��S�9�ُ؏[h_��wy^˼Ϟ�-�����>���a��AZ�䞩I�N{F��%�*����U/�/��l�����^���=�H�h���T�
�� ��Q7��Z�.(�� �WDOPƢ.�6���*�Ζ׋�ʄ9`_��_�Yz,1�x����%Cm�?��s%��d��)�=�M/T����D�p8"��4"�Tt��I��<mU�@!j;n/Ur�T��e)翻�:
�r�X�{�N7���,ƫ�W٭$���w�z���� :>�z�1L(��C���G�frм��Z�p��D�'�p��<&�y���
�9Ґa
g��6^��LS�����X9�
)��p%�h�+Ȏy�k�؛�/�W<b��$�@YҨ�^\e'�35����P�B�&����:�;�l�{C.A�#�qz��v)d�����^�=��ů̎T:N�6��o�t��F�n�0r5���&���S��E��!4�D�?ĩ�g��������os	*$��(�4[��k��ja�Y|d������4$(�Ȯ��R�忥ON�ѹ�Zbj/AU�k�L��ȒkE��^P�;nu$Ow��Z���;��ݣ�wX���#���f��w��}a��2>kM�v� W�m��r	�w~�u�a�:%��V0�����%}h��H�Xwx���1ANJץ�ݯ?�k=����{=��m/{��K�N��ɟ_����@���]9_��ʏX��_���Ky��n��`��8��[n��N6!�QM�W���� 3$�����13.L���)�F��5�G��`r�H3�IȺ?+Cʹ�y��ϼ
v��i�����E��v����@�2���j�Zu�P�'�`z�4��鯳����o�*,4�Q��P����=��:�w��T�=���q���K����樄�8�E$O������8��h�N[�`���%������s����W�	�QC?�s��H̴f!�5u�C.�L#��m?R�j��i/��<������fN�c�\��R���uq����w���}:�F{��C{����w<�ą_x{��в��da�ʟ6��~D����� &�g�"���6���¹?��ė/Y�(�o	k��X�x��U�{� ����=9����Pî@�ګ�	gb6���s/N/����maQ�8��_�Z����Ӄ��q��-tqyQ8�ǫ0|���o��`��d�\y�A�8Z$O�3J(Q��N0b�'�5��_�Ch;�b�����Hby�>\:AF��,�0;w���z�[��1���:x	�|m�χ�C��c<c�{B|#��]��_%�b����e���yYcc0K���5��#F�U(%ڬ)֬��~��F������Ｗ�����*KJ�]>��;1dWS�	��M^S�m�����ur��a�Ve�΄�a��,k��˼im���=6���<�P�SπDG#��a�ز�q��]X�����%�BAY���P�7�W��@;dE��u��7�Ց��Ht�_�� ��yϠ����F<GZ����Th5��;�b����0��/3VA�Yyj�Ǧ�(`w��#�� �����|�[m_�0]��"��P�È�&8=��� ;q���_x��Q�b�SN��Tu-����E�wE�8\ξ/O�F-�H{����;"�{��=t��,�Fk��(X,�GaƖCY�b"�j;+�Ke�_}���f��H%m��d8�ְɩ-��@U5�w�*Z�ꛦ�?��Y�q�E�I�S�)B��]��ks�il�����1Z�f�<��,���?X��۳���X՝&O�v��%T��>\�l>U4��751я���;Z��q�-!A�x5�u~��+O�y���)�Ca���߿�D>6��#�̼w��M]x�3\����ј�Ҹ7f�H	���ŭ���{(W��p��������azeMB���M�ÝYsں���O,/v�;��~4� �k�����/X#�|w|q�=!w 7s`5�`ޙ"����#��W���ت�Ư��y�L�� "`߸`gT�j���G�9���֊g���J:z��Է�`�����κ�~We_������`*ʹB�3�lvT��L��{R�݅nz%�>B��vS��O}�Yi�.gI�΁��)$�:9��/�]�!�$%�~�<��
B!`����ݸ]SQ�]	��NpQ3��g۳�������N���Z+S䰆6�'�r��lo��$j�2��Q(�%�I�d�hX���l���f�������RK˄���T_�
T��,�y��D�1#��z6�Z�Y�י�S���h��H�?'�[����8%Բ}�7��T�s<���p�#nkm���jJi��E3N��3�������H�U��(��hA�Χ��T�/�j�i��3��r�:�Tly!8Bu@�Ծ<�M��G�b�<)e"�Ct�ſ��WT�Ug��:���a�Dc�'��C��q��eْ�*Yn����Mf����f����'�L�������W�R�3�;� Ь(��i���?a洨���r��jFt�#ϴa�N��R�o�����龍�<���@�g5>w3wM��n�����Su����hNޭ�DQ���M�d%�nu�t.#�{���� ��8���홏7@��
��D$گ�-��_r?�,Z��G<�h��|�����WҨj�>L��p~e�78s�24���tӝ���}=l�gb.�̌����ɘO�c�c���5���:z�<vח�Ԑþ�rW�r��u�҈�h���&�񦵊_�4ף9��/K/��YM�z,9.1B��(�Cg?uQ�� �l7���2<�_������D�Q�)g̭��RG���.���C���V
�o����ƴt���7�Q�K_9����О:nPЉ�A����Nxҽ_5�#M���L��f�f�
Am��j�#iRc�h��6�J�6+�:��Esg��POC~���u�0H�eŜO8�p4Iu4���Ĭ�u�ߎw��Jř5�4L%������%�m�������\�a������ޚ`��`(u�}�@�ML�%\�o���v �?�Bb����mg�-���qpY�b���&�i�W�C�Q���/1�K�+W�9Ig7� ��7,�P'w����z��w=����`&�.�0���voF�����Ȥe�[�����`=ޝ�����i5�n�$S���j&�x�/�L�JzA�I�߻��zQ�ޒ*�[=����޳s7�`������o>���^}�:)�Pu��pݩ��|�C*�Y������\�:~`p"�WG������_lyP=�h#}}a:��yk�"gk�O��#�j�B޿�_Q1�w�����Ȯo��ffK�����刋K�h��&f�@G�d��Vfj"^=���>U�A��V7{dS]R���y��>�V�.���Z5UG��48ptÝ�� ��$�L�j�5|�ސ3�f�
�~.ц��awq��FGD�}���$�ܲ�o��h<�v
�l�F|��aR���l���|�'�A�D�y���(�(uu��i�������p�yW�_�9}(�O�� �nЦ/���l�k�z��6�Ŕ�NR��� B�*=�kg{�G�1X��ӾIz���",�n�~�!'�A�v}��%js�`�;F�I�v��S���G���`Y�G6��h���sC�,y)��l��R�s��Lo�>V�%���ŧ*�he5����~zE����54��H�$[��v �1n�p? ��fx��6RY��>��-��^	s�h. ufi�L����:�)��[�v��mp�����X\��#Q���ޱ���Ҵ���8�������n �1l�����f��jM�&X���al.���C�����	_w�UI�-�oai�͚OG�TGpS'��$���բ�NzZ[�*�%��}��1Uɲ�?��XF�/h���x�G���@P�`P�qL��Y7�B�G^:pi�(��qF��0C|��35��@g��}XZ;���9I��C���*ܰZ��J6�`�Äĳ����=ױ��&�bi��Dc-L\gʽ'�w���	1Fe�h���S=-���P}L��ी���Β?�x���M�a�%P"��t̸�L�/��Õdf�I�|{��`�JC�mp:�B-�ξD*a|P�~m����J��i�or]��L��;�$��p9�>��]�v�B�-|�MgSnHe5	@BB��A����ꅌ������:PD���r��g4ŏ���n��`Ӕ����NG�������7�n�=໺g(n=�_)^�T�K}�?
�/N�O/)�8��;��	NX]�@�-2*�Ij"��5B ��EJ���A���*<@�)�q:�[�Ud�^�M~*u4�'pN	��/M/�h���l�b F��ɴ8zK`�E,쇣�"�]䨨k��L4vk�6{��9HWs�Q�>�}8O��J��h��4"� ������\�@���7���%�6�9鼅�Y����R�yv|��8�
���n�,�	ER�?._�JWO�M .J�R���ݒ��2Nӵ*��Q�I�uS���U�~�ָ�"���͌�{��MQ��[>�􅳦e"��{:����a�u�M��,�S8{����ȍ)p"+ZpI>[_�1��2��`Ji��
)��4|�[䄇�_������U���0)��8Rh�O�b�3`�\��>)��r��L7��l��Zq�(�g�yCC�n�Q����J��,�� 4`�ݷ�uv�����S��\i�t5�'�s��z�5�_^uɋE*�s�.�B���&�N�Nl�T�x��:�����g��'<�J�-y���
�u/��w���yR����_JK2;��dz8r�L���eewoh�|��5
]�� �jߋڀj�1�nطx�cJ����#e�Z��^�Ua�9�E0�/^�[��-N8�������H�wG���ǒ��к���!��$%��<�p���򲪵z�]Pt�����IS�[�vf�	�v`cf��T7D����&�����_���6JE�D�'��Y�g��w}�����vv�=�LA#_��Y��F���n��Y�U
�v��J���+��%j�(Ve���p�Ő���G,<�����P�~)�v�"�ou�����j6&S��2م���%��m�$�نE�puԱo��&�p�5���	.�
?�r˼�S@��$�Aa ��Wp��<n���P�Z��=�k<��1��D{�n���;}�8�A��a���[x%K��2=��n�� ?���I���X;��4
��|�<��]�]PV��	��+8A��I�Vp�rc�ݷj��ߋ�\�6�+.+F��M.45r�A˅��j�=?Z`5��0���պ'\#�x��[���Z�˝����w�;�̚��,��3䍿qɋ�/k5<i��ar=�@|C�ێ�~�w/���^��f�]xK�S�/�#7���?H�+	0�B~�H����p7N�k�ZX���=�M�1��-I��  �X�r}��62����~��[6�Lѝ������Hӗ~��{}4��E�BAq�(�����YܑR1��Ŀ�sXק��K\t�ѝ��d�	���	[뀆���^pȇ_`BY�a��~1�ڦ�d�4N�1&�#��7���DlP}�gwg���dy�JN�=Ґ�T�7�z�_�Ȝ_�T�5��E����Kޯ9y�E;&��	lٖ�-|+s�n�D�Y��h6�V��,�����j��2o����;HLJ������Y����~2I�u�fw�A�*ГE���s�e��z�lM�PV{�YL��$c\��@�\�o5�]J`DW\�ձ�	��rH|�!��1)�}lgl�>���rN1����5����H��6^"�S�o]Q�U�/>g<xC��d�j4�i]�7��:�:7.� ��I,NMm�����Kv�#_ҟ"f�>[{����&��FE��#JU3� ��x���t�I�{7����8�W�Qo7�3�����k�=�����n�(4���m�4���Wx�F�L�?>���q"�,���Q�t��\d ֥�4�U	5��;lM�H�Ԅ�4m���#|����S�=4��dp��������(T�:�Ue���{v0��g�?..m���c<��9od_2m��Eg9�G��a
�c|#j��]���#G����P�3�ʋ�N�U�S$���]�uNb�Nv&������$�7z�9����=u�Չ��n�y�u�)�2�G|�q��d(bi'jϸ�=���¯���&�sݪ 쩆�C�Aa��P�R���1@����d��k�� �릅P�R�LC�oh��ݢ٪��J��(�����w�Ȱ��'N�NQa�&�r6���D5��tvY�cd�`�["�����
��N�RD.���]�j��.C����3�Tͺ�]�RZ����C��Շ
M�����]��R����X�M&q��S�5��	d�(�mmm�����q��rkĚ�z������
7[?�����OA7n�50=�X+,4k��B��B-a�R�Н����E �6����^�_�"��t��0��v�) h�>�T6�����*/w�AHw=Md�z�L��� ��y��q&:?����/�,�87�\V�h���sk��'���.3�w���![�����z���&��lG��Q��Ӳ�L�He�����^��M���؋��|#�`�Y���q3X�z�����Q�1�����ؾd��q����ٳӃ�ḭFC'��&g�_Sr������4>-���b=��A<g�7���,}C����O�I2:ƖX�h��L#o�噂�-�
�0�ҽA��κ�&R٬����|.l�2 &lr�U���U���&��Y�;��VqTuF+����_h�s+ia�n�S[�π�!����4�K:�g�?b��	=t1��G�mM/&��^RD�<������'%�!��;p(�j:�(Go]���z���U�W�y�u0F�%`��ǏT�l�2'pj� �,��b����&�_�>�IQ�����xd����a���-��� fV�?�	"! D�v^�?wׯ�;W�o����%�p��W�z1Z�\�.TW�3Mv���J^��#L\���v����@�?�\��}�$���eZ8���(̄
�?P@�#����s^��g��D3�.fL#�C��@�2L��O�n|z���(^_2򰡲`60s�u�O��<��z0S����夋�՝���ѐ���`M�Nl� ���H��н&�bD/�p]�2�.p��%,���
��cC�']u�rĪ�;��ie�?g�O���w���E�z��k|E��E3���];֊�|ƒ_�c�;.�+�:��D��8;�Ը0�d�m�v0�4G���������{�K�.�*[ګ3�1��k���y|=蠺������o���*C��V�3o$�N�r������1�I�+��Y禓y'�+�����a�H	\��= ���� �+Ч��Z��ī�[��)	d��s�5`���/���9���E�PH5 ���"�s<�荥�?���S��w�e�۾��>�4���@�~˄���ҏU�����7 Jx"�V�9N�zL��	��y#@Lx�@W:<�뵔۸��o��#L��Ձ�J��/e����)����yqm��Ͷ6Q'#��P�+-K���z[j5!�aJ�]��C�g���Jy	Į:�2�sB���Y��9���N�Q� ��r�0(h�z��BsO���p�YJY�z�ɧ�;8D:�(5�v�����W���:�m�ʞ�C���x�X�T1�]�»� ������c�%��Ggհ���>��Rٍ P�育�|\���]�l�Qa��-�z��}lZ�HD�R=��ZPr���m.f�OL����N�I񼘞�����av��Ia ђ9?��]��J��z�N�>J���%M}6�;V��]�0����|}�B�i3�iZ�  
���k%J���s����p��%�wy@Ռ	́yxJV]��mp��9o��������_K{(�~�=��&���<��|i#��g"���� 7?i�}@�3�F�G�B)����c.������v�&d��V�LJ Or{M~�����:4cf�x䈋K������Ը�Az���_d���3u�;c�/x@anoU5�a4��g��42w����j����%���|�ε���1-�V�J��XL���.��v�t�!a3sr6�2{�e��څC�_YP�W��f���q�VWEt$��ע+��#?X5*)$��-_K�ӗ�;^w���
�p��/M��W_�=��>W���T����\�^�]����-~ը���@�r�z���h�'�;�m�N��Db��'�@51{�SGM}e���/��j%��i<���\��{\ia�H�׼*��3\�?h��oq$?<t��|XN��\�Clo�ʈ��}�h���El�Y�8�B辱��Z�<+I�Aڢ��\�Ϭ�Dk�`��MN�{^�+o�V�������Myn|'�F�`���V�/�r�i�Z4uu����@�z�$n
i�Y��z�IVբ�hZ�?ꗵ6X�:^��iw���vztg�s��`7?��;ـX�E^��\v�i�zɋk��A�A��Kn���u
���Y}}=��~�.����g�p%a�	��w�`�Ka��CvȰ�6&On yd�����jȎ��kN|�і�|��`�W��f�cr(�2��2�J��竉[ hϥs��ƀ���&)�W
�蹟K,π��ǋL��i��ԩ�o������Ž7uۍ�/zRg;$]�|�r+��c4!6�t����H�:'s	�{~R�
A�Hx� RމOA@[]�=��5�����~{Z�-g�.C�f�y�!��O"a�;�Ik$�j2�|Q�Oq]�����<q�u0y���9I��*�U�P�&k0��:��<��!�04��>\���UT��Lj=7Sܥ���Է�|wW,q�u�C�!h��|��NP�V��3BS%�=��cŐ�,���+U�bx=}Þ��z��W�N=�?���P��N���'8�W���ҽ#�ñ=X�v�����M71����!ʭ�-���Xe����PweZ����r{0���?��.t�	uPb���>Z^ b�%�_��:��'#�-�ٴL�j��V+��?TЂ�oL�gy<��*��Y�\Ωw��O�Zt���.���w�v�����r&�0�R%�ߟ�fzk~0�9*!���&MG��$/h��)jF���6u͠^�iD�s��:=4b�񚴿;�n�"`��|>��T����cH���y�Qڼ.�!7��G���7����Ϩ�_]{HjJ%�M@�{�[�{k!4�Ǜk���� s��=]�|9oΌ8�t~��������ۂ;j�
!`�v�������+�y&f�=��:ڐ�-0-/\oI��<�/�=����_Nd�r��	����m!:#�׽��d9���7�@��Y3�[�*��=������y�� 4���>��'6��>��ORp���Nm�qh&�A�A��R����`N�����(���P����O�ƛ��9N�����jK@E����*᪯��RcA��?�e�ܞ'��ͤ*d�;<����='/#F>�[��������� tR�N�B�Y����ts���N׽�QLb�����Hm0�ٴE�����6�fwHͱ���1)�@�t�����JWh�"��#J V�8r~�X����o�qg�%|J����E��m���M���8��l1�p�/�s*'��D{j�ױt@(�<IW��ձ���L�_w�Mn1F��~"c�~�3�'����|0=��2�]�=�4\P���?n�o�wR1�t�:3��o���ET&���%��DG�G~^�B&X�TMX,'p��JM��y�c���E��c��g��yi��@�d}@���͡�()�5��)>����q*)qj����G�)�K�򇼩f%&���г�̚�zV��R�³�`�������I����{m�H���/|Zjx�K4cC�H��H�O3g�Ժ��H��!V�YS�����;*E����.n�-�� �x1QjM]��v�����u�����O�ݯ"��?i�[�^	�9�	�oZ���vy��٭�BW􍉱"A�~=!���(���5��92蝎B������F���{&Ze��:\XG�4kB��7Y4s]����mZ�2i���):Jx�y�Q��A�w�%�t�Y��z�"Q��P����E�@^�G���'�n��(��E���[pz�;��7���%�td���6�w��e�^�L�T <X<@ǽʜ�B���f�_�C�#�d����ʛ&�=�E��3��a'l���^�	���;�ܣw���V�&W��E9��Dl��k$��c��"b��O��T]�,º;������d�`�qϭ�v�)�s2����'$���%p�ܵ�8���ˆ�/#GC�|/�F��9�˟����:�F�Vo���6�Y}�ȃmEh[9�^<A��2֡	>����m<�
[�J|la�#󽟑�Il����'���@�N���M>|���=�N�쀸��i
��)��35 �!�d���:���l���P�@�J�Ѩ�U��y��W7�"�Rɨ<�d�v@}tL�@C�D�����s�5��-�͚�^M���s'��Dx+.�J���*V����^� 	�7_�`!Jj&&��0eV�>�'�;|(�N���z��l���0(����*'�p��?$�s>��d�Wӆk�}悠P�.h�~~�� p�^&�_JJD�޶C��??9�s	ll�ΜQ�c����6=��������S0���Hޏ��@C�7w�{��t�:��"/`���g����������UN<��E��B�nW���P멟��RW}������ߖ�����o�e_��4$���nU����+�d �c�a���aؙ��X«ܘ��ڣ�#�(l���m�yVj�0�(D�P��&�Wi|�T'�_��2�7�I�!�7����8�ZZnNV�NX'%#8`�RM���� @r�gW�
����4��n�+zn�ܲ�u��ɔ��>[Dv�e>6R!��w �2�ݢ�U��R��GJ�=�|"��p>ky9V?��*MΖ׏�Wm	d�.�H�u��`w><�Ъt��ٲ�Ӓj�3�"I344�	�C��,dF�nւ(���e��s�q�w��R�*:�x��<Zz��$"�����&������L�e�@�3�]z�������^��x��!mq�ɖ��������#s��[R��U�/*W��9n��7s���Y��g�y�<����e���n���"l��~ j s\�9(��Edf��Fu��EJ+��_o�_>����B�7���tz��
=���a|\����b�Z��-��l4C+`��2�q�V�߬��4Eڍ[�a�[��-��0�����0X�j����j"[�	+*&f���9E,���C�����Eu[�\j�w=�L�`͜�ÿ\��)��<[���,,,�8��&X�����������2~<�hu����C3����K��evǒ)w�?���-3�~����ډ��"*R%�'#?�m��Ղ���[�?ZT��bwe�q� �3�S����']]�u��_g+��Do�DBLz����e�.�ok:��V��_C�T�����]������$��$���nyk� M��Я�m]�I�Oͨ���%E��f>L$$��/��(�N�>�o�G2�Q'~~����p}��nt\�#g�G�7T!a��OU���_� �V�ӵutDlw1A�Z4�_�l8>e|����k��n�'�|�H�>�4L4z�6��R�}é|*���4\掳8��t���j��w��P7O�c�)�.&*��4�W5s�?�]�H���52��DWD�y��6���H��JFLVZ1����첏S���\�?��L�M�u�?h��z� W6<
,üZB�\1^�$iC��qs�
/����iߪ�,Ǯ
iGYϘ��hB��y^R|$�G/cW�D�Y[Y����O93Ⱦ��*FR�!�'pW�'
�,�Б
��=�x�#ɢoF0KZ����z���{�LI���zc�>��w_g��H�4C3��ن����I�߷�-KF�r���ɡ���a��g�[	��`�|����Avjo�gL0#-��j�r��V��#ڄ4E '�)�u�d=7V�^wOU�}w_���_�32R�x���KHv��~�׹���8�c�	�<ݨ�;Ym�tI�.���9��S����Ó�0'�eЁs�^ݻ	`�����1B�6�f�e�� j�R"C/>e�z��z��Sl���܏�Go�[Or
�V�m���H�5��Qo:��/�b�x���V��F8�1�O����{��_��Hkڟt�|�V(��,u]��+��`:f0�מ�+ �wΗt�����.���G5�ve�Z�	����ZO�u��������U,0(|v�?���F���m�(>�sxҴP�P��b�Ĺ	�:H��1X�ع�>d���&�o�l\ o��>���<�(�Ơ��2��j��׉r�8䏫�xeճZ����4ةQ	����pwF���8I1�JO9�6�*`��������]C)�v�׭1�@*������'�J*���c
�K�>F)p��t�[T���!��H]�@�F�hg���h��e�~ߦr"��ǰ�״�4Q�%�.d;�m�_H�G
��$e?� ����G��ܞ��W�����>ߵöN	�����ژG"7^��u��p�h{�<#/��}�Yֽ��Ce�D�o�X��>�If�x�2lwȉW�I�R��Tӄ�v�UC!���쒲ߥ60ݶ	�؍#�_.,��[����xk�T~��$�P�r� �:�Gʋջm1��D���``0d5�+�M e9ݿ{�h���}���P����-������S��p���^O2�S?,�91;�s�>�N,P���,P�j��cyP�LW�f��́_���h<����S�qd��z�p�]��{K>zz��o)nOz˻��v
�˸M���Ef�cSb�'�B�c�?��sn�I�}�+s�����1!-�'�����zx�pY)�3S��4��R>|���g�hҋ�Y���j���%���R�4=��1���42�h�������j^}�ޓ(�e^d�+�kO� 7G����9>�,�el�5�?ޤ��s�5gg��;,�S�Oz�*I�<�8��E�V�A��L�e�������� ������Ǔ ��i��F��i��Αx/t(��Xx; ���UTy�v�џ����7S'�]�}�ƹ���c��\������KBƷ<�����fϸF�qL����Q65����VNZ(57T޳����)hT�4^�f�*���I�6×���eۗ3��<2�;N���g �"7j�B��>�>J�<���o���tg/��RJ���F�����_W|#�G�l��m�wmE�,ꥧٔd_qU3��ͽj��K�9|T*�v��&z�{#�>E�nD$����cl�7&��n.�ux<]�%|�ԗ��'k���� ���t�r�~⹰�">I,�Ys��f��P�C��yz2o	�Nsp��T�Ѯc���D��� ���/^�6�$FJ,� T5z�}sg����x��?�z�C�od�Iр+LԹ��lko3}�ڬ���(���X��U��̸T�h���%��A�����[��jb~;KqI�e2+�C4�d�o3Hȧ�����a�h��27ێh6q�#f9��ޥ��@�B�vL��߾��l��|�ӊ���g[�,N�>8dX��Op���f��Ezȁ�M�k���ã��(?߳/_6��& ��Z���4'�0��0�w��`��E��7�ڃ�aR|�U��>r�L�.�1::&E��3?7Ac���	>�
��a�6�ëȑ��Q�hyzJ^��5����}�!Zy���
�JZ]��ʮ� �����D�#��� | =��
�V��
��mAxnN�s��Ͻ!���7ov�<`8�����z�됯�S�N`�Ŕ��!�(V�<>zz�QF{}~J�Q##�;θEEc�5Ҍn����>��mIՌ7�⊴\˧
������;V�w���נ�ќ>׃���F��U�Z�<o��\RM��$7Wk��k�O�^���h��8�9�o��&��4�0�5��ڊ�yr������0-�h�����,хf�ik[I�y������ˑ+��ϰJ���B=;=�l�c �;���a���ӈM� 3$�^=M��_��<y��H��!��r� �te��'��-a�#y�l��?a\`�Q,�/Z|��Ԕ?������<]��A�.!���ٳ�)禆�W�^�����KK���ňR{D��r
�?K�=� ��>�%E�H�_���%��y�.t��_�z�qD:�����+2@IS8ל���0Ľ���#!��A�ɖ$b;�����_w��޵�:��)�ل��I�ޙ�4�a��ݶ�K�}�Ă��rPA߆68�`2x �'>���M6Ӽ�����w���<|�c.C{Ɗ����m=!z�h�M���y(mpG����E�I�0]��{K=T1n�����~-�	��x��'�?]����2E������D�}�j���5�����]v�Y���y  �==9�|>_���3719D����I���x���c����q�6��]ύJ�G!��S@��{45Mʑ��p��Eԙ��l]ta�yl%VX��D�
\5nF\�$���`�r��<N�>���m����Ո�.��p��i��?��潼��)o�K���[�aZ{dHHX��Le�E^�6������J6��։O\]E�S%�M��|��g�ЭK��r���yϓjoFõl5�����C}���5�h�_� ��v|�W�9�OX%��_?�t��Y���j<zMG���	weD#�5����G��E��u�8Jy�Կ�,x.WM�ڇԨҝ��������:�� ޡv��Y�=_�V�A�>0��)%B����io	�6��m>@��PD�N]5���A$=� ��;��>%a�Xp�<������?����g3�\�f�+�C�f¤�.�Į�Q{���<6��T���Ч���:;�q1�	��$d��.ێ�*c�㹛�MWТ�Lۧ'}�Y7OY�\��9��������[��H�'�B_��l~�,��:f�^a��t�]�&�������#�_���/�jX��J�^YP0]���;?�����]��+�wc�k���~?�"Y�2--/�Ck��s�pFxn��1c�"z
���K���KMy��x��aY��d*�Q��\�5��4�����#˴�v�H�C���6	9�A�#�ύp]�53I��V����Ƒ�O���(� ��ov����d����Y��u��g���O�/�y	*�(�5��i!�W|�κ���䪰��΅��P�N5�.��+�D+b�o���f0s�4=ܓ����Kռ�l��q�A�I���ح��d�Q�,�0Q�����{�BÓnȪI#���L�����i�d���s��l7 `F�AdH�W�͑p�ٛU�;��MFIDD��k��
ھ}V�����n��۞i2�ߙ=¡��j�J2�ho�Ϣ�w�b���OL|D^�wk��_�]��z�M=6���Vm�M�e�W¦�z2x�P(�&�'��x/g\������v'�?^<��1����̅������w�����~����ͥP̂�=����� ��mp��(��{v��Ӛh%J{[{�@��xk���./�d_���u��k���A�~�Zds��|ծ��`/Q��̌=�X+�ӯxW.�ջ��#�O�r7^��?�޾O:(���`;oX��P?� ���2^��S�Mvw�z�N4���	��*鏌LAf�k�?UǞ��1�gC��Y�+����W�����X�)N��E�P<E�歒?�� ��$�[!@���n�o��S�rO��0�SR?��ٴ�3ᰊ�����ި�ޛ�7���QC�A�� �G	�f���Ѵg����S)_�R�ϷW�j��� �ɦ�1uFұ�B}���\���Z5���3�H.�B��d��e�O#߻�/x�_/� �b3uj94@z��Pt�{�{%	��P�eQmKL.��|��u<�P�7��_6�����ZQo������;ͳ�
0���5?���+�p�\��]+nP��y"v_���Op�}���Z�*������HhJ��>���"�l ����!����޿�lc�u�Y*���}�셈Bd_�w�dK1�}�C�2!�Z�>��u�����>����=���<�23�>�u�s]���u����z��s$=w}�I�?���0�YN�C�e8�ι�לA<�L�	G0�en�Uc#P�-�:@�{�f���-b#�d~�x;����h���n�;����j	に��dS���J'�-��(���(���R����؍�f8�xR���tt7���
Л�G��2l�:���L\�I����S!2���b9M�oe�
۲�X�Ht�Z�W9V���!t���l۸(
DyӪ�Ǎ��)D�T�vaYdE���c�[NQ�t��;d�>n�_��;�Վ�h�T`	}���s��<��>E�.
�O~D���A/��;�A^��������8��4\�ơ[5�?�QC��RP/mE���IJ�)�U_�}{�X�X�绤����&.��I.	�������̀�G��R���Z.�I�{�Z��kr,��z83D8H��e2�����6tm�mt�=Ɗ�Ŵ,\�eϝ7~?UL΃F���+��]��<G�Fn�/�&��ݏ��<�ƒ>yo���ֻͩ�i>���V	IJ���#�N�xQV� -��G8b���>����B�J��j�8����
�<I��W��;~��E��꧶�z�4j4�D�_�P������K�،v�)N�ؼ(�ٓ�=���O���Iq��3���P�a�،u��;e<�т�C�M\p��9���i����R=}+�z\��\���$بs��i����OI�����r�d
��vlN����a�u:����k��2�8t�"<�2ni\�uP����n	3z��qlŰ��<|���IH�	9(\FH���Qk�Vx� j>^-ߺ�y>:%8�ж�Zؐ��A'S��)��l[}�t�x�ݵQv:m��Q3C�Q��-�?,�=�eiQ1l�c���y1"i�����]a���gB�/��5,�/tŸ́��7�Q>pde|7Yv�������0���f�]0py����q�Ǆ�׊�[ oAi�U�@f�/�UL<�;0�+�_-��=`C��4���t(� 20���+�	�~)�lE�ߎ�I���P̖���s$����O6�T��5�&�̡���ci�zů����:8�9��ԶF<��:�]i��;��@͏ڶG�!��))��3X��?�b��������i딫<-B4�{o�S4�� �ڎF���S��X�$�.,&�.��f�ey��� ɗ�&KpY�^���cDHm\�[�z��F{Hi\^�
�;�#�6�#�s#��<���`�A�fRvS"Z �p�bb�P@�����|���H����X�WܷH��/�ai���mL5�.p�@��=��ڦ��F�uc�Q�xp�7�l��������x ucr�);�|��;��У�[�q#�9́�k��G�H�L@�Ɖ���)%��0�#r���qj�����m�/���r�ɍ�}AlyBӁ(PCs�偑��J���Y��+���L�P��/K$VV]���BM:*���@�_��|�Z5W����hڥ�I?�_�o�r�L��cB���"N��<�E�09�W������ӯ)6������x�]���+�^$,�r���G��Yك�B��z�{-�cVV�l3j9@}���%��<-�"��^��h�(���ϕ�[�N#�<S�_�����Z�X5��N��c�<vwMr����Hd/�d>��m�������5��2=��ޒތ5�G�8�����>�l�La�`#p��a����>�A���81E~>�p�/�[. �_��I��5�3�#
�Yl`TH�Ss��v�`�`6ɧ�wW~d�v����A�v��`��e��ƍ�n��1l���	:��x-�3}��|��g��u�2�������\�X�8��V�3�PDg���Q�3Z`������	��]�*��mB|�ٙ��T���0�~�lQ!�lr���O##��_ȇ�Ɛ[��X��]6����;z�Y\P%qx@���/�'������:���/��a�v�`����ء��݀�^D��[>+98J�]E����Wl)������>�;׿��j97�E����d�n���]�a��WT���B�O�]��f���w�85��诚��W*:��d�qN�����N�58����G���&����
{Hp�j�7�T�Ђ�zp����a�֎Q�X㝎�����[���(~q���,1%]V������3� �00ܢr����!�4²��ſj��ٖ\k�&x�Aͥ�{��:���)�X��Q`�9S�6+
��O���ך�������ϛ���|	!����� 1?�M������b6ZN3�K�������q-���1fh�h�|�J:ի�1&<l�~v��
yED.;_¾��v�uh���a�U,��~��)+��S�@�}��Rq����|�'XK<��h2.����g���-�����o�.�#�1qʧ�M�y�	�u�B�3S��\`�G��k�H�3�V#���׸�KQ�I�4=��복�����9��o��Z�M�v͝�@�7��V����t	i�z qv>���#�h����G�����@���:����"��8�?�O�v?��3���������$4Y'�0P�-�Rgt]ȉ��h]���a�/�� Z��P���k+��=��1���� K�`u��pG�NN=�r@���{�5w0dP&�`�L�6��%++��'�C�x�{�l�A!. �Y�V��Ň�cN�2H�ڹIp��:�ɑr� �k)��g�X�<G�*dR�?��+����Xs��v���=4�1��v?R�.��[߇�<]}�$X
rqø��D{� �OG�ʭ_a:{^�Q�f蕔ȑ��@]��g(���b3M��\�!�5Ż�0��b�wJ�x���	����ٸT���l�r��lB�G!'�V�M'+�{�`�<�R�f��O���I$�u�#3q0�uu�`3~�ܟT#^��.�����x스�L�
�*Va���=^"�;s��jV��5��`v�*��FD�����i�(����&��\����܂Ӄ[�˩�(�0�{���2I���ɱd@�}��Śܑ;|T�B,ܼ
睦��<k��&��HBx32w(�򛺟������]�7��=�@�#9%�#�E���z4`��e�a�������.�x3��@�T�f+D��ֳ���ԁH���̉;��8t� ���E���V�:�H����Rj�5�p��]�>�6�\�/J,x��D��w��٥�q��˻B�ө�~�o�)�+ݶ��f�գ�6W��8�yH��:}9VM�=�iy�w���$39�LJF���Gx+E�Yo���F�i��f���g��@�XѨ��8Tw������1o�+��S� EXҢ&Tx�V�9R�&A<uOz���[��Ξ�?��]>{�V���<�d�g��ҥ=��Ӻ���Fy:���t�l�� �{�yP;ƴ�^XQ\nY^1iFY~�];���p���EP��Xb�Q����	��p���~�G��s��D7����Y���`�H�#M�A�76	)���W�+C[5���*�_�AVT��STǭ<dF��{��m�n�[Br�0�v%X��poMӲ�����Ϣ<��/��Q���K(b�����
]Z�V�q�oc����-/�G���`�#a�� 9\�2���QZ#�)*f��֤����v��#��[���tn*hET��\��Oׯl("��~m+g7�g��	+���0~P��&��ma���eVW�>de��'&$,�X��1l7���9�<Զ�*t��*�����PȜga�����		��d��=��h��['Z�ݐ/�Q���_]�s;[%�s[�����=����:����-V�/�<�yI,��8鳘OV�<�K+�:F9V�ɏ��?��o���=\��|%s�yvv]T֜�5�)]��z�`��*Z�+�}oib9�Q6��O��[,2�}���1�d�������e{O��2�4��EG5I�&�5x��KcsAy��%���ڎn�*ml�H)x����݀F�S5�"�X6$���~��ϐWC�!�ǃ�lU��P���Y�S�Rp�ݹ�OY��>>uv
k��S�k����f�э�8�����[��"�����^i�ӓ�XZFD�/..�3�=�N�j��|��r����4�:GOO߲"���������q�RR�x�9��Q��fd$ˏ'��S�S�f�C��f���Eɑ�<����Cn���M��t�⚌���#��mв@[3z���.V��l�C��1�?�Ya���#aл��AHV�3�(&�愅�Ggu�,/PGA�G���Nzs���E�|��t�&t.p��փ����ZmQK?NP�'���OYP�υe�
�'7)�)4�V>wfEMĐ5D`V	�k����� �24=,��LLW��+,�(�Ei�Ӣ�_Q,?0�'���t�k{���~��ؓ���Mb����eP@]U�lև]����K�_���$�s5ڊ��K��]��fS"��(�ݹ��]�	�+\�u�5�0q�iC8"ϰ4��Q� ,:�ص	�׸��pbu�y�N�P���X	T��t}�᪡�_-}Y�AR��k�U6h��B��L����uz�!ݪ+��Uשy�6%)�Q�~�����R�?
��(�������|�kT�8-M���l��}��E�9?�n�QO��ʪ�<��|}>����ܰ�"�����ӵF���e�h9vM��H��P��������a�[��4G�ݦ��]*f;��}�{�y�.u_Te��Aߧ�l"h4�
^l�1��D�U��&����B�	�4�m���w�Z�׿mШ�Ȃy˯�3�N���w�7.����!yR\�}����?Ōz�ܔ��V(���q�{������JOkA������&?O�Pf��h����e�Z�,�aĘ2���ަ�[��_=�_o��|я�Ft� ����׿�;���a�b�Y��Fb��D�wU�Tc>tٴG�
4�fUT���Z;��)X�ż��SvT!#����L��M?�
�9G֏Ԡ��3}�w�L�KD�p�G�ݎ-�'`�P�*N�0Ю!�NҠG��>z����y"�"�2�.�p�rs�mL��>�t��]18����74d�cK��g���^�\$-[�����Ծr�J���IW{9���Tr��QC������f�@�WJun{�\���ڇ�8�
�J�t����|0,�<����P���+a�`�n�TT��.J��M'�'��k
�s��E�g3�~�m*fGIN6Xj.�����DnX�.$ِf�2��hG�:G%���V;���}yI��Ax�R㬶+ou�\c�z��0��<�1�/C�d�4"i�^Y_�{�jI?��y����^ $��mβ�@0��1Zx/J	�T�y�p(ɫ��9{��+?J.����<�YxV���&V����� �ӟ=�M��0�~ZD�
o�+�}��F�R��^�Nz�gwuu�.'d@yn�b#�w�+���L�#�Yj�W�x��
���'���D�=ƆS��S�%����%�	q/T�NG��-���c5�8��j!�l_wwV$F+�W�cb����?�<:8�^1]� y��QD�����9QC�59a��dGS�':�������M��ۘ�O,T@��;t��"Þ��W	�SiI���A�x��D��ʈ���=I���=o5$/*�0�%1�jMe�?n+�	!����G#h�E����S�ʡ{��nK�������j�l1�!�n"h����������n8(�p�w~ո��>��k9��lD��6�t���'�"W?�Wr(��~p��'
�ϔ)G�˗
�?��n�������+ A�h��X(��"���6y�I==Z���vWF����˯m�\Y9.H�o]}�a+�M�{t�&`��SKk�aU�������6�����C;zb��_45ͩx��D��!5��s��9���1ޚ5�G��*� !GFg��|�|2��<����w�y�pa�A��m�,i��?�@5�,WVd]ݽ��F�uTA>��ֲ����c���gh[�gƞ�ݰ#ҙ}z�4o*�4�K�HK`���2�G�0�n
��&����9��U	�âp2/8�]�,����k\��k��q{>m���T�z�p���a���o;��-̻ZZ٠9�� ���O+�Y�J��^��:�U3�.Jקu�I쉋O�C9Z�s䲢v�Cx8��X�|�6���f/"K����X&e�q+����h����5x�aC	��W��/��^�ǹ1GG;Y�o[(�#�]
q��ҌX��X�&�fv4�S{�*�=R(x����OG �P;T�����;0P��k��W,����cإ�~�����~��<�GY��_ߏ�\.k|a���J.��G��>�C4�p��'��.~)�����8G�XcyK��;7�}u��۪V�W���j����_z6��td�<J��_N�~�wB��'{�d.5��a���͛J�LV�ZW�o|y�����ϥ���T&T��hq���;���yO�r�\��B&p���>��Ӌ�|�: w�r�r��~�RW���{�	rhvzT_=�j2�f�c����ʅ�h
��C<U�e9O#fo�Kz
�me�����w=�H69 T	]��>�3Afk����ѱ:��KCC�^����M���Zf��I���L"����l9������-�ú�{V��_�:Ĉ�痿\_�n�͛Co�	^���._H,���|���k�!���\cp�@ǅ�I�P1m�Ds&�FiE�m�{��7�w �ܵ=�Tk��o����1Y_ޏ2eR��P-��Ւ}���A�@e�ȡ��A�ͮ��d�gPb�P�z�o����$��;���\���f^pd�@�޳&n7!�)�}��w#gnhn�ǰ	��}죨���l����R��kf��Ѣː�蔲��{ɣ����:tA��/�OE�$�A�[�h#��X�r�N�{���q����cLe1G���/�}3�����V���&n���7�!�6���(�c��p�0�p��.�T Pw���Ll�P����"P����_��;�_W�-���ug"�tއ��B��S3�.fFe�.��@Qa��B�?�"�+�u�Je'M���q��cWi�k'<M��Y[�����K벓|T*5o�bEJ�#WË>�%��.����FJ����|ݳ�OO=���h]^*P���>�����g�s��ϒu9j�M�c�lS#Qt�ׯ )�~�4�蔾�D_�̀I0\M����L~E>�,³ˮ7l��5�s+;��9f���<7M��x1���frn��pR+HT�9?����'\5p*�&"�� ;��[�[���>X�-B|#����s��!S1^^�	��JׂEϯQ�sf�K-� �Ѷ�yZ4YP�czFV�>�AR}Z^�
�X�����V�`�t&��x=*{sI�i����J�c�d?�Mjh~<���E�TN<t��¶�{%fwV���mĬ��̗��F��M\W�݄���\�u��?deqZ���h�s�����'L�^�v��'�+d�0�(�i�٫����gF�m-��z���g�	X�Z9`z�γh�2ջ�7�\+�ܾ�:����}�������>�P������W'.o��ʑ
�Ƿ���
�����#p���ö�c&J����D�����N���|m��<LQ51]F�`-��)�&�:l��}��.v�k�*U.s�i�U~���������j=��l�g�ۋLuբ�`3iǜ���o�o��>Ѣ>�9"ⓖ@p�k����Gm�àM�ة�����\']�� 4>�1��}�{��b��g��ĕ�1�=����h��4C�<�_m�	����QQ]U�K�a��â��/X�yu�.�W�l	Z�L]aoPAJr{�1y:�ON��)J�v��kD¥ �tg���֙k���)]?�f�S�Q�v��=�z�y�Q�`Ӯr��qr���&�9n.x�G�
�P?3I�vQ*��G�9!ق0SY@]�˪"tt��{�Ə�)���b�.&��Lt�o����g[���;�"��B����Ձ��ń/��X��f+�7���ѡ��>{�T�"�l��{����b�G�|������%)�J�����No�F؛�[�fAJ��v��4ǲ�dYrM{?Mf	�Qx:Ê<����L�d^ ���q�p�5nx���4l�w���ev2jk�6	�y1���|X�gkr��	O�[A1�+��HO�s9��o�
�B��P4e�[!23}��5|�����	��<�q�"��{���4��g��4�Ch��|6�vǺ��7���������ʀ=("��m31#N�ī1m�r��%f���搂]�`��ʕo�Ve�[��~[0+c�C����Mr��_�pz����3.���L.BL��@ĳeٞ��&�,�u �I�Oǆ���ig��_n����|�nތ&�@���F��Z�R���&e��|(�k:��p�T��'��X�rl�PVE�sU���Q�
�6� k���_~�bywM��5s����v�'yq�ӟ�1i�vcq{�������Ů���.�TtmN��U�������=uqb��<�^W*]�"��f��2I>�Z����8o��(1.k9р�D6巷Hw\�
��g6�S($���2J�U�2��PR:n��iD��J��oUTMB�(ɲ�ʬ��Oo�{�}x��>�D�h,c|Y�it�����"��jv�Ĝ�x�|xCB5��j�606�<�9~a�&�g�HքG���,�G�%�[v���l=�&�'7���O����Ҟ�9��R˶�#0�@�X�#�{����}�w1�B�_h\i��J��8�9.ɇ�bZ����fCe0�M��c圼���Hi1��fl��":����""�r���5��Lj���9S��輹��rT}�v�ւFG�2&:C�B��p����2�����XoLGY4�VVV~Sg9�����n�uXʃD^Ͱ�^�x�=f����퀆SQCuƘ�d��7u�X�M��}J��5�4f��ş+\*N$yY�h���J�vWW�JM�v�Q����ojFL������ �t����s��ono6$�8���s�m{��������(+�5=���ԸL�i��8�?��H���Wx�MJI�>߇������8<��y�7��!��pNE=1�본� ����\A�W���S#l���A�T����q�a�-�Ǉ�b�lp�V4��������F�+�g��m"�|�����l<j�é��c[�6������WQH�C�?'dK���E�Kr��"d����r5l��UyT$�g����ï��@e�a�+�ի5OF0J���1K�g�{rO����n>,��HP7��t���C7c�ǁBzͶY�u��$�Z����~�я�\��ʑ�g�Q�g��xh�W~�h�w{�Zk�����	��}���~�������r�r�֎�QL�\��!��ӑ`��#���7���n���n R-����-���G�[�)3��i̟%�!��B�����W�y�U�fa���E?P�K|7��6�Ωm�6���5xl�[�-�H:��mEƆ�N^����J�Q��m-�W�9�%m�����D�u���VY7��-%�,JZg�O��éشJËU�mԼK���⿯�U�ѫĎ/m�q*���\�ϜbSL�`}A�p##ǛJ�Ε�-�m��F�,�C������E�%�s�.���W�=h���� �f;q[�+:��΃��Q��@#�*T���y_�pvgwq�Cݱ �hD�l��Bd���e:�/3���1A'wM,���^DFZ!X5�Kn�~�{Qh�e8xk�=�%�{ʁ�4��o�e�x��������"㫅�F)�9�VI�nw����ſuT\�����j�e�W$��GN,��6���?�D��ˮ��Ν�d	�U�e��x ���a�����R���w�M�O:x��䕂��X�[T\
o 
&~w�bn9F�/�,�=�~���JI�P�k�����sc!�D�1P�xM�,6�q�&<��gW][47���<�8#aW5�"���1��M{f��VL�����P��.�%�Aޜ`�)�j���m_\^�t�o�8���)��uA&�k4�E>�W0	��[L��=ۜ�l?���8(XxOz�>�<'����������a�`��c�I]��X�Z<�7�M�����TWᱹDWYI)��@N���}�-�j�����$a�z�D=g�>'@g�,��2��j�$�E�.���R�PRe��ܐ�͏��v�k���]WzL���tjV��1��,�`�@8G��=��Q���ׇQyK��9���ֳ)����!\��ti45�_�#'��{�A5���^8«`o�O�D��u&��z�|��ےY����t��;3�_�E(��r*�j.�K����R��$���G(�G��+޺�컉�wl�v?R�<��[�Xbn.[�s�D��S��(�-�i��F���(�gZc��o�c����擻��fuj�f;rAE�lcbA��(f�n�l"�Vy���5Ʌ&�de�ʷ)~��qun�@�X��)/��:j$�N��By�&75�v�{��s�S7�a}��ޓ����6~		���9�/���Q�/,ƴt�@��2��E'Њ{ob����5{��.]R-�ό���"�[�}��DluY��ļ��l'N�R���S*7�ʈ����I��T��Q<��������e���;�t(���ܺD��]B|1s�<��K�}Eks�΀R��.4���H����u5Prխ�ږ7�I/�r�|�S��d�wR�#O邼Á�QC�^Fz%Zn���׺�].kL0�v-���U��'S:L9����*�<1o,����O�����E`��fԊA���ܜ���ً���H�e�}o�@�6>
���v�a���2�@Z.� m:�
�O�!:�I��&�bb�A_�2'O�ψE�V[�dҒ��t��x�<'�oTH�X�?��ױ��E�D����%Jԝ�,D�*��ƀ�ڛ�����@ۂ�l@�6�c	�I�ED
(��l�i�7/j�Y�!��J��Z�,�;txay�Q� ݑ��G��j�OƉ���JZ�a�F�-�1���Q+�7:��65�fN���N �����m�!�z���K��Y�f���t֟���
�~w��e�)�<9'�y3�HA-�{p��B
�'!�����I�����Zi � J�9�iM�-e��T�H�|��T /b/JPlߎ87�A����dT�t��\�D�9�80ഴ�p_�t^ȯ����Sf�a� �}���XR�ƣ]LH�c�[���ce/ڹj�w�%T�a����%R�s4ɪ�/�,�YI'C�4�!@ݞ��	���6��P�{����+�w�)q�?�!
��ļ�ڌ^�3:w�=4�"��yr�0�����]�5���u2ף
�9���ƴ�� ~*f�v��^����K�
�]u�"
�"0,Ԧ�^���(�שu�xT�j[dwjb�J�AFr�
T���������^�B�(�/b|�c�/���㦖*ێ�G(T���Ң�3l�'99���"8��wۣG��j^5sR%����Ke�h�V�~;�_;s{a���L�I1�`��Y,0�F�a��u^XL�R
����ߡ�*�O�!�D�z�B>%� ݸ�X��A�*H����a����l)�#}��\�*V�O;y�󻭔b��ܘ���6R`ض�Y0��Eq�v:�
��T~m�V��W��T������Sa]O�u �*}/�KL��2�ë���&5��DE΃�p	fw���_�g�ٷ�8��~d�@��з���3}/��j��o��)���`	��*�����"���+o����	=�
�t��\�a����Y/��_���I�8��?:��&�r��*��e����"0�y�;G��l��:^U�W�T�eb��6ga�j5N?>ФX�L�r��찑�`g��x@f�O�[#�����@�Rh�`�
$�YQ�)���H4X��&߁�_��o�g�ሻ��Z�/�}ۮe:'�CG�T�5ȿ�RqK�׬\��J���Gj�栰�P=�p��$4w�
�|)��d+������l���LZ���D^	!��Vq�G"�lxxx9���}ܩ�f�k�3�Xd��'���	p0��l꿜�g�'l���x,��C��ZD��w.Jf�{?��C��#=���xjH ;���g�"ѧ�>���4&T��姗�Յg^��Ԝ�S��̆�mՒ�f��#�c+�"�t�m��r�T��Ō�6���e@}ԫ^u�]��،�vno~��G�k�5�^�0~-`�Z��-��t�����C��R��jM��kIm]����.y����i�:&�� �U?$c���Y��fE��8���g����{si�u'U�%3߬��>/pMi���xp�>^86q�� 7���]gC0u&%f���_3.e����D�ˬ���k]�s�l�Xx��Dg0r����m&�6�/.��h���XBF�iӽ����$��Z�����@�\-�5=�pc�)\P ��@k��p����r(�O����O'����W�#���z��}8b�d{�{zL��Y����n1�t����(_��MLl�ǝ����W��_\�:M����ɾ�@S�ry���*񒶻�?�d[\��/�@7�b��\�&!��ã=a"���8(�<�-�ʉ"L���D�yY0Tau5�(�d�95t��������~��⩆���x��7@�B�U�miX�D�/��*B�C��坎>N;I����E h>���AF_��o>���=�"l�O5�Dub�B1Zk�ғ�@��Ϯ0��=E�FV<xbnAZ�^�ྲ��i8���<V-��`���1����ɧ����F..Q.�����g�
����6���30C�c;��'T����"���M>�m;DP����KV�p�qD�1�8^�H�92\������b��e���؞OD �>��x�4t��q�����wO��o;|�c�w6�w�^�M]����E2���n��,.��y�I�T�E�ĩQ�b*iQ
pdcm*�گs��.�U\FwXҡ�j%�DHuKO,�;�M���`O���|r��� �Yĥe���������:�$��}L�X��^n������b]J�Q���o@w{����)N8x8%��kQ�3�ڊ^�%w85�4��r��
Zo��>���g�r���J�p_�rvj�(��{쇞�c�;�ww;�s?t�Ɣ�!G�nm����}�b���e���i(Jn_����p��������~sL
c���'9.����_��\�/܋���A���8W��/��s궫>dzrܤ$!��~�;'<;",��`O���v��|
�����Ԙk���ì@��@C�٥ ���a		`�����.��a�I��W�����6��*m�Tՠ՟:��h�}�_p��I#�h�[ݜ�K���c���1��|���N�(M��e�aE��'��D$���/��e*u%�E>�l�*Yq�ˬ��/�o�G#"�?>���g�g��i�Q���y���Β�Yݳ�2S�怃-z8� �% ��yb��M�ⱼpjv��[.03x1������čY��ǆ"G�t4��e��Q�c�@��6��j�F#R�TH����0L55���_ݔ�(����4�u���co����=��u���~�~��|���߃�I��#�@�q��
8bNT�ӜG��.9��/�ni�����#|�L�o�l`��&�*��5����C�=�w?fc���M�//o�1��?d\�Af�.�1l7^UVUY��ͫB��ѣ�w�֣y�7��s7�B��<��AVD��RĦ�_p�Q�V<��qJ8afd�WR�.�ȃ��Uw���r^��X��`��; �����9匞r�l�}��璞��j.{nLe���9εǼ����WòTe��a`@���ǩ��� K/ r���6�ĉD�ƈ�9E(Վ���|r�D��8����7��2kd�e��9o�2��Z�����A[�w+n�V�߿	]"D	��h�_b�����m)l�l�07&}�כ��-e�
$��ȑ���D��1-JD�@��P���'�|i�~1S��p�k$C��1�w�#h�F�M��[����=���VR�Q�_��ۅ���c?h��Vgh���L�]�m�����ѱQa�Y��D�� ��b[���H�/�R!�Z���PV�4ڐuS<�JY���9���}Q���l�$�K;>"�ۂ��IZ���H5=���q�#�T�d�(������bm�v"�@'��՟�πx?�ly�U;�IQQ԰�9�g
@���bA�ٸ;*����}���"} 
1��YX���6.1�2����6~��wO�X.������9�[��@�q�s����g��ֹ1�x��4���ׯz4�K�ʘ;��k�3%��qw,��%��tS���2S��ɑ���0�HBIӒ��j�{%V%`7�܍mt��8��+��������Q6��=(DY7����-�h~�����b���w��~d�M�c����dJ����4(��e�]���k�b۠<|������\ꞟ=����[��3^+q���22?�o߾-����R�f꽳6TQ%��w{�X����ğ�]R�뗰>S��#�����_����XA�	��	���{�������_�^#������~��Is	h]�k~wI;-)Ӂ�U��{���������@)����������Txk&�c*�q����W����i8E���Qts��ׂN z\ޓ�R�w�UU��c؅��Bt��8���y���<��S��胐�]�m��̗��U�����{�W����d�G���x�C��a�yja>�ɵ���]�OV���N�du�w�w����
u��&�8��7���@����|��V@��S�y k�����oA�d��Sɐ \^wFc�A�
�Ss��஗�ì��2�y��Xbu��.\������(����3�1���np�^D��v����:&}���w��]��y*��τ:u5�
E]Xpj�`��
V��,�ܴ���VץP����%�s�����V�Q}4�kg��[�ݙ�:?J��A5�I�p0 ��S�g�g�Jl�5�`���6V�bϴf`K�kD*v��Z����?h���_�0��s�17l�Oߖ��ݗ�I�|E�B�j�@�ֹ�<#�L/Ҷc`��c�<��V�{"G���W�pd�09R�ʧ]��.S0tƠnD%��ڡ���m�Ŗ?q��z�ɱ֛�$���3���b�}�����ʉxh�5�1����ᝏ��C��O��p�H�s�	^�<�S��H_�)��N�.Do�~��`�X�Q��lD�~ QA����"�y��Kf������FWH�7�&-�q�q�{y�ses)��R�c/�)���C9�����L~���122�N��J}���������_�m��(ҁ�Y��a�DMoh~8������`�c6�<���ݒ���gu���l�A�\pw�E�JSg�0MfRv���H�}���ʏ �	���w�h�p�6�,ib`hx��Ux!��U|7�����{^�bͨ���o��8�:Umxχ+,��;�*�)���`eB�4��c��s��}�87��8�/��5lѠ��}󳼁�v�m0R��*��V��
��SZN�Z�.0�-��Pg��7��*M�Nm�:�N^j�h�a�
騍���n���D���j����|���i����Ƈ���O����woi�칅�p��6]�F��Q��"3/$y�[��;'a�{8�l{g���y,sGS�9��AM=�<��@<�u_еU��]�mQ0R�&���^��֐z|�����Ͽ^��ښ�����X;3� %�����v��~W�:!����b�i���r4���Ǟ�~ �)i�zĘ#���X��_��O3�aEb#�&me��ЗP�c�6~�t9�z6t��Ь��!4�z��R4s$�r�4P����y�v\.�.�2���w�A&�
�.��
Kț�r�1l�71\�~����:}?A���2�%��r��'-�.������<-�"5��(%����k�]�|��T��p�mG-�a�1�7پz�y��r~�ާ���iw��Ջ�׌����x�x�Ռ&hjD�eⳮ�9��z�W�2���
����4��(5U�������\ǸP�����Z�L���*�~��ɐ�|
d���ɾC�vC	c|o��V�P!�Ǉ�6s ����F@�C����6�y������F�,���`�������3��݊�ۿ���j����<�<��)���WkS��=�NX��FC-+�x����U�ʮ�B+t������#�;h��{�b�{?�59`�oM��k[;����sJ����V�\���4�jWA/�.�׹ׁ����۱�B�}$��r����) ��v�����7Ǥ�m�8|������k �	-7�C������!t�Ma:o����V/.=�3݂,��78�-/�{)�>{���-t)6��t��x�X�=ꧬsÌ�M�\s��L�]�u$sB��x3�b(�U���=:FZ������M%��CE�mj~�;�ܡ�;��C	qS��'bo/��\[���N����(k����h���m�'Ll�A/�̾8���铖��X$��CqaK�﹐��_un|~��1�K�*���Y%�=��&0�c������4���;�N=��^�|�����4�㾤���8�1 j�A-���-F)��� ��8p�ߒ�������[`^01�*z]��Q��q���E��U�&
��x oTj�k��ЩC�z���ӟ��Q�ހ��A�A��]ЪȢL\2p�^n�9ܠ�sG�8Rs=vG�2��.��{C�V�n�����uZI�.��ǩd�T�@�ϓC���O->e�somڜy��F#�x��5%�<�g�_ x}��p�$�a�c��=ӷѶ0��H��q���Oʚ�QJ�ݾ���>����ӓ��E�?J-���`u�9�R�� �����K�=��{O��?��<����,�-[��PB���(���bɖ%B�}ʾ�%�u,EDٷ���U���:C~�L�������?�לs��u�^������u�ɵ�^���c�s�"ڙ���@��z����1�b�����}<�hpm�u�����ʌ}�����y�u�l�Akc������I=�v*���@�x�W8�Ѱ���Ɂb��ط	u�Ԍ��Cl��5��htN�����<p�4��x�,<O�,1�&q�'<���(6%�jU؎*ZXju0B��'�~�{����ܫ\�ߛ��.?��Ͻ�Њ������"�S�}�'	�Vaߒ�	FG�xƛ�`\�k��Zx�"�t�����%M����N�X����1�>Z�:;��M#�
^cZ��	m�A��x�X�kUv�A̼�p��2{#
Q�Fq��Y�9L=�g��6��mOК�}i��6���V"��Ȣ��^;�xC�eи�BxM-mV	�j����9���U�D6�lpM rꧩ1���C^x����@`"LCx�#(omy�sZc��Dpr��C�q��NC������*���L�"��V6�/��R&K4n��}�U�	����7��o�u-�'Oh}D!D拎J��0O�	ݒ�������W�!\;�'�T��㎨:���-W,\·��n� ��d	9A:����π_�{xS4Վ��&lW <�Ωt�K�H��s�\�U�#X���D��R��+��P��:-A���xDs�p�iQu��Af-�����]�l���0���ӳ��d��w;<a�7WJ�X�,'i%��ʔ�[kX���M�ptQ=u���ܢ���I666��)�2B��D�d��G��v���(�e3L2<��\���c;�]�hL2�İ&���=XN�p}k5���|J���y8xv��ٌj�+��;���T%�֒���~l�.��W<p2,��[j��;����q���{iM�INIkw�H������e�t+CR��8^zQ�,�Z�U` c}6�!]���pN3�?*�ktI�����NF!�M�U~��B�]������4�Pq�Kd�C���d�bbP�{ub;|����Q��;HڰƎ��S?
1���-�K��%�yV������rz'����H]b}~~��1�Ȯ�J�R,�&%Q<z�B���m�?I���g+���f�Hm���^��:5�)��
�wl|���KkA ��r�7�yҖ,�܃@�)]y:�����κ��[��n-���鷳/� 1�f�e_�J��o��j��Q�B͔��՝��K 霐�tۇ~�q~�&DO���}խ(h��+����Ԭ��x��0�f{jf�,��,�kM'������^�EC��=�>��ߗ����ʪ����+�����sR�\,H|��;:p�V���v�:�a*$�p��e"C\p��˳�.�,�z�����^�qh�Y+/�dnyH� v����*\Z��e~���{���1,U���{���̀�+ �^�q�E�H�<#M�H����.��2C_��'�K�Y�c��"���YlX'�3xE�e]r���g�	'��7�Ŀ"��|i;���J�ޟ��.؆KW�מ�5�[�c�{�?�'�Ġ���>0j%�*ȳ�T�J<�:v��ruǯI���5����_X�҉�%���[K6�}˩/I׺���mmE&H%��9*r}Ev1�:��0�[{��� g��wp��k��v	4_�>u����|^��3mt*�#�AtI��|�ָG�,���'�$���.X4���XS���aͣI�D��z�b�~4P��[mZu(�=|�! �Y�vw��W�\�{�! ��7/�ɻ�S�\!i��/����v���S�A�ʃ����e�A�)x�'s~Y�9�/�U�5l�aM�U����ڦ(��̈Lu��_����D~�z��Z�_ACc������F��9/dU�>�V|�a���b�4���߂�L4���~��#��^ir��/Ӫ`i,�	��I��`�9��n%ְ��J[My�cA�|��v~;�td�uu�>z��=��&�r�U�̽��FP���d��wL�%����鼱|!e-m�Pwp8ݑ��/�٫(aVu����s�^x����,�˴2D��J��`�1�cߟ�`/�|V�c�('o�R�͊N�B��)��2򚷃�}�u�Y����PЄ�S	{.\0��J������C���l��f���i`>q3=�zw��.5sߤ��ϣNa�e�,2�F������W�+���[G��!�<jk��3�da���&S�Ѩ"����}�;H�q@w�\�ar-�����,0��_�-R�}�F�l����е|���c�S�44��R<��gm�t��~��1�����1�A���e��g��:��PK�<�co�9�?��B.X?�#,x�C��{j�)\D����ix��;	�=իm{'�`LA5#yG�ī���;h����~�q-y=q�8}��@K����ӯ��]pwډ��53l�O�TD��ӌ��o��K�57&-?�H���F�k瀧)���$��D2���1�O�U:����xIJf��W��6��s4��\�Sm�.qd8��ϗS���i�ܓ�x�Q( I�ӆ�&�5�p��|�1�۳+
�?4�T�'w�b���W_ ��\=k�:�8��vR%B�������[�)����z�RL����+_8n>�l��bk\�w���
��0��+��#O���h�����ZB�
�f�ᩭ�?�v������J������L��ю��O��/mg�N��M�pP���f��ŷn��n��뎖ode��OU���Z��#��Z���Z��HS4��o�������Ҥ���p$�"����+��W3Q��-�8�f��}���K�Έc«�� �����U�e�S?g�I���*���)!��0�eW��7�G�v�3�&���=��;ۛtB���'`�8t�N��ճ)uGq�y_b*���!��� ��-1����)O�O4���=o���>�1!����iXh�3��q4T�V���#�;�t�#���B3��RI�m=8�k�q�����Zʠ��$aּZ�Jg{Ev�hma��J��o�]!
��g~�� ���vLWh�'leSzj�X~!�"
����?�K%�ŚzW��d�j���f\�ʞ�;�-�_Qk��r������Szۍ���� �E]fP�i&�N�E�E��TM�����.�:�m�[��pZ���K���)@6��}%|������&����W�|&�6�忩h�9��%�;�ӛp���0���TY�Y9����B��G�j��G� 6��D�W�d�p����L�¬
.��lm� ���X~D}��F��k]�&B;�<&�s�.�wvgQ���U�͹��d��;O�����k�с�s��>b�d�G�du�I߉�Oӈ�0�İU��U��%�����O�����x�[_#y�.��{�Z��u
�	*�+��0:%�g���+rw]<�o�$95�Ӹ��D��zֹdݲ�]T1�*�ݜ#9�H���N�o��y˞s��\v�\����i�A��o���РB��ڗ���֥��$��I��h~��;o�x���C���![�8��309:G�����b�ףO�g՚�G���w���Q��b:�@k*�4�Tp��9��)��٩Sf^�]e����a��40�����[��a��{���� �]h��_�{-�9tX�v��g�Zm9Y�b1r�%���Ã4��Y,ߤ�W�x��^�(e���D� �bv+� 
K��]��v�[�đ!�d��}�2��+)��C���Ѳ�U�Ę��l<��X��]ZX�@VG>��]7��c�U'.}�A�D��˜t!i����ѵ�o���B��m�o����5]�>G�o)F��M�(�#R����1���ެL����&|�7�k)��}V�?��k,PNFE�]�o���ݷ�~Ztr��(�>;����>��a�Qm��k�t�Z�CM�26�
u--��'K��N�Gߞ�NvK߷v�Z� �";W�={���:�)� ��� �3{����9΄߯6�o(���}�$|#��l��qH(Z`Q��9cbj|�]��YJ�"�[I���#Ϝ�ŗC^����Ԑ��`�I!��TfXa���t�y'�<^ZL� f�C'di����OIp�H&`�P�L�p/K�Rj ��,d���2�1!l�<+L�#��jJ?�zL�7��0��e룥�y�%6��p1Гv��+�@_�O�{�X������,�㚞���3���R�`�VIk�d�65��Ο��}F59���[��0���3�e"�_�crN��*��xp�9Ԫ|}o�g��Ӵh��b	$�	�G��U����
����RI��
�����w�R�	q�����`���w >G�`c՘a����"c�؟c�T4=�U7���	-�D�M<�eЮ�X�����؅]0æߗ$Rq�q��?x}ƖU�*�'̇��������IB�)�.?��C�|�v�Wا���FC!�ew �@b��j��г��$R�ĲZv�@b��������x,���J\Nn'��PS�*��P�^��+�g�7���7��)<?�o=R����w�� ���wE����;���<��5�˨&"r~|�k�]ܠ@?#>�S�zWL����O�~�����,�ѵ�uǏɄ"�O����`��@�y�t(	����.�
	 �d��S��:E�8�9�m%_�,�i*�>j�s`��N|��>���D�#+�O�g�wu����� �+�<�nt���v�����h(Yj�}���ɾ��~�Y[0����qa޽���n*i=��~-p����Vʞ�V�G���Y��B>Y�$c*�PoLM?[Q�LC��H2zP[�GZ�4k������Ц���)Ca�T���\�&�5SR<�&~J�MHF�����݉%.��(�H���"�$�o�f�>@y�����u��Ф��X�|%�'����x�,���8}��x����o`����=�J;�2�D��C���B��J:��T	=ܝ'ME�z�Y�>$Îv��S�Ⱥ�O9�b;���x�����\!�4�����af1]<%#�� *�Pd��tE�a;/=�=kJ��O2Z9�fH~��8�Ǆ���A8��U|�rt��q��#0c?����HI�uԪ��I�,aL�_脞�'??�[1��7ʧ������ϕ�g�)hP�a��u.[|"����]��b����[�����:1|�e�\�O�-�7[�n�ׇ�Y��/T������nU���ڀu�d�����r��MW�{�5���:.`�E�8
��b��dT��6'�])��� �J/ncp$��ˑ%�֨�#�7
���6>�����I��m��n�����3��V Qb��~��f/�Fd��R���B""w
��ǽ���3%(1��^՞��aUn�#��s��
��Q�_$����%���<��w�PԹm��t���]W���]����ʦi�߉�K�y5�-U1�ufH~t�g��^�����oɺ�b\	\o%��N�ӈ}�a������)Fv�,M}^8�y�Wӏ�����'���e��s{T��D��T�#��g����sJ�����; ߯V*sX�����L�ԯ��,����P`������\i��ٛ/����z����k$�s2̣��^�wN6�� 9����>Љ�f��~vuщ��ff�	ۡ9c	������#�¼�y���ȝ����Qs�g������kt^�4����K��DA=:m���BFy�3AM.}y@4��\a��9ɨF�j���y!Ձ�����REKR�+	��h�RU�ZB�XU�o�3��.o=Rx��e��
�+^)f��q,���tXQ}�N���w��O��	�|%��i�+�0^4~੨��V��C�F�AE�z�Dq�}c����Ө��vn&t��?�Z̀�?�����߂�2�\�<
ގA��({R�9���Hsz�.���>y��5a����*��e�����>--�<�'c.���!�b5��}k?/u�[6z�x���Ży=A�LƼ�BaQ��I��~D�z��� �=��!I����a6$"N�ބ&�Q�u����ECw�0�>@�����^\�u�9�ʖ,\����	�����ܡ��s����ngE���a�xtR�t��E�i�{pi ?c;��`-n#�/���C0�@4�H�l1!�(���}��MPM�ge��R����W�x6�ʛ��,��]�����\�}�]UVv �C,�o���� c�}IsA^np�C��;��/��i{}~I���1��vBy&Oɛ�A("�E��^e������v��@��3�F뽋w�Ā2d�*M�^�B�	�����{��VP+�WK�M�<�̬���ƕ�d:���d�b8Țy�p)f��]�[�C;�ۑ�{�[G�'n��-�@��&I6eI����'w�(��߲��j�	P���l�&�P;´����`�e@E���H��B�lN?Ñ� ����\�!	ƃk���Heߥ��3Ƃ*�,&C�[�0,�.���%��=���ܳ9�n��|���vV��l��Ʌױ�߾K�a��r~��Φ58��ځ�ARw���-Bd���%��.�s$pɰ`���zL��kD�bq�S�RM����9 �1�'T�Vh�*�}���Y��_a�����:06\�
��2 'Hn��v��}�?	�tHo����)�T8mݷڎF^�Y��G��E�1է.1�jͺ���{�S.��M@�3&GL���b�f��}�oK?��N�O���mf[�JRרI��='e^Ӵ�1U��.VO?h!]+��v�ᙊ!H���7k��W'�n884�zZq�3���O�9��O�gU�E����x��]�6~��i�G� c��ME*����"�\$�����@�g���y�JpF�q�T��p�5l�%�0�E��0j�q:�c0�s;6�B��m��q�r��97�u�/:įk�}!�U������a���0�^�t�?5�ڞ5|�!�S=E�Q�ꄸAU�껵n؄�
A�n��U���*-,rx��r�� S{̈́B����N�u��D�cp����2 ��9��cJ��	��`Df��� �zTz�(f���"��Uc����
oO���L�YwV�p���i�3\0m���Qvx<ϰu����ffcs��^��[�\8j.#v󵒫e��̛� �西���w< �����|�����*u�#������0�C@%�8����=Om;�9�Y=!YY6ͤ��;���B"��0R�V���͆ �����m� ��������M����/l��׌�Ѱ��	b��dp�h�$�~�̰�t^d��?��}7_\����	�NH@���J?�n�L�v=�����$S}�w?oC?���B�������]�Ӈ��~!"�</s���jaw�g@�7b�^��;k�h*m;���f����T"������E64��eT ��З8�M��9��G���QT�� �U�h���M@Dè�Bw������E��f�Qd�E�:����%�Y.��~)�xq�c�Ol��1��Zi����"pef�U�)B��B�R���a^�A��,*:��?(3����_�=yZ��k��
+�qO����;��ǰ�Ö���>����@NԆIz�y�J�)��/�[�įh��(���-�m��
�v���\�W��=֓\�WHY�U�y�o��̌�6޶*�l��:+*�6�{NZ�S� ���P��}D'|����d�H��o�nc!�-1�"�m'.��p��G%Җ�J��@�K�2��еC(D1�� N\EnԨ#a�e��o�EE�Їo�ċ���lF�'~��Fh�k��-�,0��a�&��s�'#�w���ۼY�]�W��(Bn߁(�R�l��
}�<����)x�ܧ�s�}Ƒ��}SAx{bku�&#N���8�A*��$�B�o�A��	����������	�{$��NReb8�'�����}��E�Z�@yi���"O��~L�o�z�;�g灗�P�{)��3;�a��2-$۵��������J�y}{{�W�Q`*�B5$���0���x�m�H�����v6��0i�vݪ|q��)�w(_"N�隷�}ў�"b���� ��u�qFX�����ɖfް��L��tӌ���T 5��o�L&pdg~'��� hT_L3R��s@m�#XO������W���i
�NP:%��z�l�{z����j�������,a����kP��
�!���7o�T�#r�H���쭕j矌 �G�f��o��w�*ސ�#x�G���s4�`h|]�[�3y^pM�]�/�I���<�_R�%7쐄���V��1�����~,r�t��5��_�0*a�K��=<��nh����ޏ����	�Yk~!�{K� ����b����S1e���Í�v��y�_�{�C�d��V^%G��@���9H`ztVV�i����ǣ���ѯ��飑*GH n9���ܬ:�	��2ֲw����y�6�$�h !3v��Jr����x���S�o_��lYX���{;�ⴓ�H��;黑��~?����w��ѣY��� /\�7'�]�v��W��~�%�asp��dKB��$�'YG
 �==�ym��ǏU<�F�x��+��]�P����mE^�_�ʬ[+�5j׸<���d�X.H(�SG\{;`�vr�P6S�����������eZ�C�w�V� ����c�k��]�,��,�s�N�������tou��M�+xq��g���c2�zo��O�/�i�8��k)gcch7�E���v�����;�a���SC}�Oh�ML�bǲ/��!Ƈ�;�5ȋ{�i!�O��xoES}�E/"*������[=��N�E���(�C�|�,��i`<^�n��&�f�j�0�,�}j��t6];$>P�Ya�y���?��pڝ_�^5�����^6�sL�f�<2y	��4�9����+���Ơ��ױ�����a�W�5�&��~ �;�Q�a�¨K�-�V"c<�ւ>���b:u�"M��ƠO"����~�ĩ9וÃ��
�y���!>��_���Z�߯��)Dן�+���Ϟ�l�9��=��f5��% �=�M�r6�|ғ�<����&��'CՋ��.bj��b|��H P�H��`�v�~>����.���m g.���U���jn�|��R�乳��L.t�K�)��_�v
�ŏ{��1�ݰ��kj�
��qH�sX�@�p�i	m��!ƉBT=�b���=Gh�ѿ��O�<+v�&���C�8X��� <���}gմ8'��>��7ۣ�z�X�z��� ~>mh�#��z�Xbk����u�\�D$�A��Ỹ�ٗ]�tm��ɂ�T�^0P�w�c�zgT������b��D���r�8�u�h@�1$���weg���:��X9���[72����7���qyD2�	���V��qW�\�dU�禡ga^$�XWS���&_��K�|v��Ġ���%�5����$"a�p Ѐ_�CcG���1>�.U����r��X�B����9�<EE��l�־!��Sé��Җ�+o�9{�#Df�#��q�����E��'?ޙp�L`�L��r��k��dJ+�.��rI(�"����+��������	�πtW�Z/�s���_����I\v��H"6�(��V�[^'Ҙ_�`�Ӕ�����~{.��2o���P|ګ�'�1��f_����:j"!^�a��J�y}���;[r�{k�#ͻ�U�� N3���w)���rd�O/e4G㹈=�0� s�s�����Db���@�7Z��нrD��84'i�jC���Su�[Dc��O�q� �٣����}5Ë툴yɵ��(���
���i�����}Z����A��A��B��i�u��R��_��fh>%C����b����������
M[Dm�����e  �Bo�+g��a��-�EÏ�Q<�������g
�%KL�2�A�����yf�F�#@Wn\3�K��?���Z6��V\�X����v�M���B���ŷ�j Nl���i�c�:Ț{��#���k���W@��w�)����֒�@�9�mN�Xnn�1�(��s��3��ftې3�VT��$#`�ݸ	��D(
z�؊n�в2��N��0�����v 8�C|Y�P�I��{G]�O���9èS�����Xa��f\ z��~�HF?��iR"�FA5?�����V�~��C("q����yugBԼ�h�#����d�֖@��j���#�� ű�6u�v4��º#����w��eM m��3v !�&:Kr���~�[�>��x��V���&'_6�p{����,�y�!�8py��t��4�*�y��И	����bZU�D�1��÷��ğ����4�Zb�;��L��
*	)�4ZI�΀�3�q�553��;�b"��8(�`N��[���Q�-]V#K���T�i�E�\�Z��&�Cng^B�4^N��-i�f�}�� �E�D^�����`��<��G"����+L?5|��V�����[��Z�@�hu+'y��.��4}�,�%x6��q��O*�f�l�G�wo�b/H� ��}�@;��y%N��3ga���r�)G`0��(vb�H�r����*]J$�J=F�y��J�HA������Ġv�쳸�CLy����mnz��l`僈ߡzl�<,1o�Cvwv~��*Jz���h�L�8���$r������͟[R}��,J�ð�Ĳ�W2��*�\�7�MJt)���e��t����:��?�Ԩ8dE!�|�$kUI�3c?Z	с��W�H��F�2秢zXZ�3u;�Y|�3�iq�o��ģ���i���9�@5h:-!wp��vJI�`O�s�V�A�f(��;���C��Md�$��?�9^6ZG�_�Luf�6�H}�w�W �?�rӯ����"��S�D!k��s`t'-��ǽS����}�R�}5g�4�ɳ�g#�_6ś+A"��M�����8�F?��8��
A�&�֏ww1ʀm��Ξ�()�%ʩK"���jBQ��>,�23\0���9M�$�#��)������fT�?�/���GX�vh�ƻ�@2�LX����B� 
���`��%�G1p{|�сC�¾��f�춲S��|�Đ�����~C�,H�r+��}��	��!������C%�
S1�3�fX�
NR����`�(��6��	��Yw��[@�Z꒠��+KgP��t�����RF!����������@�����`�r@wC�;u@q\�9��<�	������p��i�H;*� ��6��i���x>U���R�K����ci4�7!A��`�8���.��e�tL
���g�!�i�0��VM�����{�4��H��۬lE������]����2�ـΛԆ�����/����Ёk+��.z����d����#��R��IS�Zٙ$��[��y�q�k�ގ�.��| ^_�{���S��q��v,���M]��]r��L����~�h��
i��y3Np�m�0�H�R���ԝ���U�DǮ�U����-OӚ���[�{^yQ�
<P�iwZ��X�I�֝;��s���)h�̊��I`�x�yY0;D�>�Mq� 7�ԃ����������|GW�kv2�~((��e�U�8�P�Ӌ�Ja�V��1J>ʻ��aHy��٧߃Ci�?�Y?(S�����۬��_}.8%�o���Gؼ�C:��Z�T~�D?�U�Ö].^V��#�N�?��թy�2s	��{������{��k�ö��<��z�筎J�/�Y�U}�(ZE!��I��^`m�	e������BW�m�\��&��Y�t6.K4wo<�R�~�����`�lw�bi�H�I�U>l����D,)22��iKO�w��ғH>_g;��sK��FT%��^�(h��*���Q|��.�v���h�sU!~�x��=Wy�t�82���9����_�����6*���5N�r�'��@w����y�p���yu���PI^w�g�c`�\�����v��o�go�j�ț�hx��T7u;%c�#t���9���)�3���?L9���m񲞘d���fL,�������Vzu ��0,�6s��������-�����K�$}�$�G�?�/zu�惹�Ox^�Q"R�{Պ�.5����]����W�)���#��&�����y�"0��>�4�U����|�y��{�n��ԭ[�7R���9���uU,0�A:��I##�9�m�2�8���}���8��8�t�۸����2���S�K?Kmv*��
�-�,W#������od���z�n=yr�o�w��n����u~�ܫ��v&��n�V/��]�Y�E��3aU�͒��'�R�9�s]��+��5�§��'�Qo���[E%a@J�LOI	W򞋼�ÁuV�A�&CT�,���+���kФd���Uw��c-�y+&F]�����d�����K�o�_�k|��c"B^�|���<���ʖF%q42������i�����R�L�_<���j��H|�B��{]�2#�FpE��I�?9�ad����i?�lQ��~�m�3��f+*���B��x'?�$ӏ�8|��d*J�7��ΝTO�k�U7S�%+��Q�[m�Hr�P��rFF!ho s��I]������Cցd)�KO�O<��f�x���N|�01��K<�K���?��ĩ(�r�6LR�B%ЉR���Q�8�Z�󖾦�xޜV���~��QYDӿK���t��$��N��c[H����Ͻʋ��ة��2��9-� v\��M��>����%ᡸ}���h�o�R=�N�-(�f���O�rsO�7�i7��zMm.���7Z��WN��K�(_�,
�����;aq���F7]L:��s�Jg����yiF�$	4�����`�����؂dF��xd]�M�Ư�Ö1��!C9���B+�:*�$@
噖w\3���mu����B� q�=����� �ׅS��2��[0褹�N�����Q�p�pr�OqW|)k����\ �]b�ⵥ�ל���q�N?J�&����k���Y."P���1��K��SO���m���� =,3�o"M'��.���k���@2%��P�� ߦ����{�w+m����B��/��R�W�n		�&��Q�RB�ـ����j���}oEA�j��y7�>+V�O���nV�-�x7�p�Q��p����9�Z[OΜ�HȮ(O7���ڭ��W�w�/�]	aG���|�Z�M� �s_��'6 ��`�]h���
��N
ܝ}�K*R���l� �&����Jn@*}�F�X���vĺiW|,?1R�����s=4$%�e���M+tIp<
i���M��s�[GדY�Fѫi�q8~�&�z���њ�Y�ry���b#�qC���a��%����)�D��Н�Z���R����L�թO_]��i��!�b�x�y��-�Hp]�}���J��٫h7��i=~�!h�4D�ԕ�����~��`�V̇O��]Pg���r��`�7o6��{1#�0��&o�ع���F����/%]�")Yk �=ܾJRR����d{�-zA���
���T�u�:���D~�D6Y��A�ݺE=�O�dCAp#��E�#-��hb���S<CuI�~����y��V?$E� �x����)_ϖ��:[��~v����Bx�0�эs�w��< �N�p$2o�*����-+,,�	=�4Zm^�5k�6?�Q��]\q
ATn�.��i+A�'ԑl�g��?4jK'� ���B���]�����g���f�́����w"��͍����1�DJ@�S ّ��#?gA�a2�w���Ënʣ6����v�����Ƞ����P� ��Ȕ���`��^K����=HZ}�^������2JO�}$"�s�o�瀖��|�q�c��]��]�	���N����]pk�U��><R�_A8�H]��ٌgM�ρI����CP�2���I� ��Y�[
�q���dC�,q=�ш��0�~��k6m�d(�+�i�O4���0뙲vt/�-��?�ξ�[��G���M'�ǩ�E��C� �}�7g�O$t6����[�
Y<�?&T���{���q؄�=�7l����;)�����c���'o��k]\8��NyK( Ԥ�gQ{�tS�_eV�T��I�p �~KO��!��弉��F�s��7���]*2�}���
 7�m~W��M���@xU�2<��)M���<�hq+BԮ�fط���Y?]F�������W3�81�����a�D�K��(�ucH���ƐEfX�*��7�h��B=��0Ba�}E���^�m�wBQ�$��	[d�������ca;��!.����|���_�A�g��L �� S4a�m�}�~0�Q]�=0ӔM��p�+��=@���3P�a���+�A��N�Y��V(P	_�̉D�8%'���x��{<���c��� %�C�n���ʹ����Q�cX���2 !�� F[�
�~�������'��\U<��l��
�l��Kʺ(�k��U�r�I�D�И�j�@�� �Qx5@�y�n���E���tb�	�dT�O� ��LI�Im�я��1���~���10V.���5�y��H��������I6#+v�g���"1��o���Ű���jX=[=���V_*�DG��ۏG�p�����6@�	Q~����r9�e4�삍:����;/�=�����@gW���Jm5���O�@�=���E
�0� .��τP1>�ƛݎ��Q���>���7�A�},�ܽ��~@kV�u����j�udҳ���o��j�oהּ��,���&9��%��|�r!��Y$���U]`�6�L�EړR�L?لv�@G�W6U�EB�+��;�S�a7���P��$##Z1r�Y����$3�����ua^���tm�gA�%V�"?�3��ӆϿ)5��'�v~�7�#A.�p<P�~��ekM��S+#�(2�~>d^�Z����o�g�>2��A�\�U�C0(0�������&N(�F�g3�]�Aw"A>����*er�w�Zݗ�@�Y�_�G%����q�vv*OFwێ��z#5(ﬠǰ�c7ca�Uv���|K3��d,α�ϟ��#Q���0��"c@��gѻk'�`�䴲����z-��VW�p1�o����Qt��]��?��_ށ�2�>�=9J�s=���:Ϣ_≠1=I�	]�Fn1�^v�Yr���I���r1@��k=Q�% �Gk����H�h���>nG"b�8�>O�'�0�O���@f4A��EY�p+�|�H�����)Ӫ6�>�A��#)U���'GەHb�w� ��"��Lg_~T"�$�]oeC}��s�7�m���ǀYF�el&���{k���Сxo�Sw���Ɨc�#<�(��PV�L��U����1?����<��=��	�sZ��-̏�����������[і<�ؕ�ˊ�bX<��ŵdeeG8���f�9Q(n+��5�=��5�=����?m�K{��㔡���)E<������MxE@��q��G{U:����q��EU����*��m@9&o��v�;�)6�毩z�ٙ�aC(5��a�7(�B�Yڢ���^#�۠B��l�I�A��2U�������?N��Ov����6#'�@b`�9{\���q�2�V�<�uґp�� ����[�߽e&�N*��X��@A{9�I�ʎ#��Ys��3��V�b.��������e�?���֙��Lz%Hs@ug�v}_�&�3r�p \�Q�a���j�N|�ա";���J�����6l(�͗i���q8�$>YrݗS#<��aT�w
D��<G#.��Vv��dB�*���
���	��lCꊡ�~
����ٛx֜�&�z�k�Ŝ�6ߟ.�nx<�fs����s#��_e�'ɨ�_3s�q>����k9	(6w�DIE���/X��m\� �M�aneP"��O�pO�SJz�q>{X��������������٢�t��N���E:���A�G/4�����[x�QH� /�r��6��G����o���UYA��/�G+�!_	�W(��c5��y!d"���g��eɌB|�3^��4�����PZ������|�/o��t��i�R}2�%+�Aq���Y�7(�6Q�s��r_�����;��)�l�H���:
���\�������Ke�'����=�
�P���:u�D��4�� �k��9���$�ԕj�`�,y��t�;�V�p��Cf�Y׻΋n��S�>Yb���˶���nȑ�XNë�R�8b
��z�<ǻ�>n�-�;�kŵM(ꔞ*�鈈�c���a;���yi��'.z���W�(����o7^%t+q��G"�Vn~7(���ᦜU"o�<)�J~e3�p<
<D�Ut�����q�\ǻ��[C+�X�̒��)P����
���-���t��d|@:�N��~�� y�L�����`6��ИT�YM�H���L��wj���a�a��hh�,��Ä1��e�m�s���IOZ9�WJJڳg�����h;q��U<���r%j�3i^�m�q�lQ�^o�ɢ�&�9����W+���h~�b1��޻;���vOj�X���a�0�#'5�T�<����ۤ@ <(P�w-~�L~�àސ}r�A/|�\Ǭ�3HH"6�8-����%��������fA��]��`U�\8	X(��ДaP4�*��s�c�I}��HiC��P��\��?���c���ѧD�o��p n�E�U=�Е�#e[8���c��;���k
/2\�Ѷ����%?���t��Չ(����_�ݎ�g9��3���o�}�]�����iL��h.'��x��d��c{����O�����6�n'�;h(#���`b�6-��'��bX��-�Co�X`r��1��v������OU��&[B�����\���Qy�������O�!I���Y	� �;���]�S��S�Fe)��E�����	~Et;-Sjff澯�Hh�6�{^M��U*Ku�\�>k�ۀT"o����7��*���/�})!��%��2-֘�!${B�}(� Q�K���f�f0�lIek,ٙ�dh�C�����������y��r^�s�s����0�H�b*zii:.��ݭ�a�s[)N3UYϲF���c��_�G���7_@W��3���찓��ѹbގ��DO
�"���w���:�=p��6WF�,�]�*�s��09JY���eUO|s�`U���}z�����1p�w��.5��u}�P���Z�~�5������ۿ�~V�5��+�'���q����f�������̯�Z�\��;^n���\k"e�qG2$���[������r�4�~�bBi{����@�\������j��C�s�,Z9�k�˘�Xj�b΋hH	���5�9���Q��x�(]�ژ�%slg��7�[֕�ra��]jU	x=�<ѬhZq����Es����o0���U���˫��)ƨc��NU �WO��q~�v� )&B�:�[�����7�L�W�<'9W�)�8y�f�k��;޵�^�x9�s���aq�1Ro$ް�;�}�-)��N�l~V��Nr����<���w������)9�O��Jz�g����i؎Ы�;���'��4��~2�i���M�t�R��ǎ��xdS��׮�G>���G<6�DGl_��n����3Z֖�7I{��]����E+�2O��m�-����Z��ǽ2M���/���D&U��R����0��e�Ks޹�dw�tjZ�����qu1K����䮬�Щ`�It�wp�>�GŚ�Ϡϧ�x(��[���Q�JJ��R��y�*�u������N�m�V�$*��ڌ�G���V��ѩe��� �	�`O^)n�J�M���'/�Զ����U>\$��*�a��y�.�_Mx��37�U�p���������h��W���s�Ԡ��9��P߰�,K�ĉ(+�onO���O�]kc��'���لs��6]�S>߽[�	�::ܫ���L�q��4\Dd��c�Ԛ�y�Ǵ4�z�u�t����uf,�u�S@0�0�uRC�E9���I�nd����g�_M��NZ�[� ߴ���0^0<<�,q�	V�g�9]�abz�f�;�1���E���8?�� K}0����CZC�����p�[앁�'�׿*[|F==BQU�7:.��'���sDw���I=ߏ�6�������>7�wX՝Ù�;#ex H�+=��7"rz��x����c�HO�L,L0	�n2��fk���W�U·&�z�a n����D����2�eϭ��w����j�aQi�Xk}W����F��`3�h=��MA�$z�ޭ]$��8O�#��ə���QV�A��6�4�]*��In�f E[�9�J�HC/���S�Lj�a���O�d�5)u�B�
�(ws���O�ߩ�w�uxV��bد�t�D8�v]"s�Qyt��S����G��ğh��S{�����2��F>4,"�̤�_��x�����_�Sao&U��u'jV0Z&�q��i��+�ƿ ۙx&�~��##,�5p��:ώ�zAr�X���	+��Dep{u
Qi��Gv	����4m��_H����(��ˑ��,0�U�<�PO+�532�aU�Zē�UUU<gT��9.X�*�w�ؓY��<����H)��*!��-p���:C/�o��Itj�7Nsn�_����j�}�`ǝ�6��s�� R�I��x���\0�IrA���t�y�PILMΚTvD��Sv���9��iuL�C��V ���ۋ�&@�E�d&�#��W��^�v"(�s��5�~)���*E�A����1�s� ��O�}Хa�u�uaovZ�o��� Kʊ��P���;��vz��c�9��M���uR��<�]Nj�6�g6�xw�������v'sΆ�������d�����j'AL���F��]�@�t�)�V�2F!B ��|
x.{F��A�̴_GSe�/O���846����f:��-v���̓��M�J26h�#�[�4�B,�����%�z�J�e2�M���=����(�Rdy -{��Z_���5*��J�����쀮��
�X��[vgb�q�I}����HT�&4ʻ~����P�y~���#���b�}�SzJL^�^�ǉ���\��:� �����x���ѫ����<e|��!=��3�|�/��A>��om������Ox�<K��R��4#v�ȕ7�,��_�>��c���H!t�:�\��E-�aW�oml�v(.fj@/��A��B+
�E,�H/G�9�۞�wt�(~s�$�'��ȗ_�H
�.��`vw��k[�?0����!%;b�l�Ë!��V�n�IW���ȋ��{�Ҵ��w��BB�.��M��	�NV���϶�_o]}�9�_�îWUT:Jn�:�o�R&��D��H���lH8״��T?��׌���g�!_	IiedZ�K���OYS�"�C+�Ҳ57W���6�������/,�x����j����Kn��G#�Vy^��9���͞^���:I��[9z��f��C�~��Wi���<-�m�#����5/��2�^yя��'�w�ڬ9�����(� 7+D:]��{�J�:�h��Ó�%ϩ���˙��($Ғ�4�T��[21K5��r��J,��ߙ�"A�_<ͭ9aD��
�.�]�:^��^3|�Kp�M��F|>_��f�w��{����u��h6�8�����z�z�iވ�
�c���
!���z��֏��Y<{M�v���q�D�R�{�^���n?.�t��Z����e�˛�`��sX��w-==���@���8��r��LՊ.���L��2����B��Yt>�q�WG�c�61FOO}f��+�М�cO޺�`��X�v���|���V�m�d�'�m�X�@�(e�ǯE�i�_v)�Bh߯~g�K�� ]�ءg78���t����r�VK��ɡW�iy��S���E�6���S,؉����x����3�A��h��^&����z`
�<66�c����un�?/9��A~�$ �T�_�W�ў��N§p{3�����e���t)⠟(��TT5P��)"���w4|���S�c>�a{�9�NJ��ގ��N����=��v�vE��Y��
o�-8�Qh�Q�ѻ��/�E���[���8.܎�[��5�;8Ϥf�1Yo��t�����n)�Qq��R����22'�-�/�B�)��x��d-��6Q[�7������eY^�bCuu�]��^ݍ7=b���Ĉ�=���f�gڬ�@�cj��{	T��&[#s����3�������x�@G�N���G�����(<���)�i��Y@���j8�M��F_���������Q���������:�}���,	H�g�1�iɠ����e�����6&�]O���Z��O
�w/geG�́A�S_�E��ѵ�:}j��_��.<C��ǝ�U��2���Â�)&MC�Q��=�v����
>d<Y>QW�&���)o���5��me�?k+�Z|�:'�g.�>ŵ�;������7VIJ`5�:ל oy?=yUij����㮡���SDj���5ݢ(����*z]{͈����E�:_T�}F�9�\�0��
:�mh�v�mgz��Ȭ$���޻�7����oB����W3���I��P�������0e�c�V�(}�>��
)4�C=C�㲃	NӚ/���9?�ۨ���?����!�kZL�v?�1����J��v���)_��7Ƭeg9�֔9�Q�9<����ņӜ�[__w�D3�}�L��Q�y�v�EĔ��A)�mhh8�o��	[���=�'r0FJ�+"��Ǡ�}bbb5�s��J>�Ĭ�'���]u�x@�^>Tz���%�[VBr��zv�_ьLh�	�Ii]�w�����酴��W�2���c���(cGY|H�݀eh<6+/�*��#�i�X7�WX�������ɣ���5'��J\`<3��%J�����1~�@z��ݻ�
kv��NnF���fwg'��g$Ġ'c���7�����+���r[�`���qE���,�n��J��i��r�!/e%y�E�O+l���0S�����V�a���߿�z��6��QS�z�K����v�s�X4��v?�����^��l�)v��aJ��R�:�ִ��+D�~�)�8�JZ���V���I��#���@i_�5�cAF�/��$$�BB�B��]��=g��r�����"��D�OJ#Ln�f��1)��P��1�?V+3-�wo�E��kL;����`�l������SӾ�w������ �y��T��MAi��yqֶ�r3�c��=9$I���1�N���iH��"7��U6��>�p����-dT[�l���NS���g�j�9:�	4|���ϓQo
𱜔�YchC�����#XTYTVWlbGG�,�\�`���Q����S��'��(�,���ˁ��o����R��o�Qy��@ ��N��A��8�=zPx�h�=���
G�2z�y�����?��̀���"^�P&�5߾?ddC���r!n����xóB�6�`�__�0�^�WZҩAz�n|��p����f�W��h��%�m����d���X���b:X���*���
K�V4��E��fB%8�@x�4[��J`ȭ&�aʛ�ȓR�w*C6Vܖ�b���Z\�;Q֘���V�=�L�jqs�Cz5�8q_�:�6��앬�`r�ԓ�F��S8�gQ�C_�s,�/�'�~�9��:��:;Z�}ІC�\u� ���D���//�ڌ��=���"��K�,�"������a�}�~+`�K�I���;NS����d/yB�aO�(YQ4�k/�| �y�m7�EKxBC��J�W�@�Fo<�!���@���vJ�;i�o�\-����p�R4�)� 3t ,8ސ�.�{�v��2�d������/ޞK��ۇ�`����e�.��d@�G�%��;P,E�*dP[�}�%p �@v�����i3�v-툈�Jb��t脂�Y^��p��Sy����3��c�a[����@��q�����rAZ�d���0��>�@>MLpkٚ=ܱ7o
p?1�AL�<Nb��Q&��V�uYr���Y��ԣ�g��	��� f���ķ���X�����I%oܣs�7c�Tw.�A���r
Q���.Z�����Nzw�e ^����gO�����&��YDA@^�E�@/�Fs��u����8x~�""��B�%^0�&��
Lȍ�����~���%i� �=D���� _#՗��G�,�},o^QN.��*��/����+~���G�~͢!��i��irC5�`CѐXT����)�B��w<��=u�W���z�r�Ԁ�#U�
�3��QN͟�A�o~��*����L����'�"y�/َ� HZ<���j!���x�����WQ������'_2��m��=S3E�+2D��?�~{��p�?��Me��:��y��k�&8�����FS�Qs�@��$n��(���&`���8�*TI֠�̀�"!]xɟ>���Y~ k��Zf�;��i%M��n[,���s����9�]�%W�"쟴m�y�2����#7�{�W�7ɗ�H���"�]������L(���@�?1Y�>��B��.���Mf�I~ki���z�q9�7:����l��L���'ك�5��">33t�d��g�"��K�q��T��c*���h��x�`�*��71��7r�����{�l
������޳4ż�;�V�=x{T���$�%��5�-��<�F%d.����'&�p���oz����V�$̊���5&���(�0��"�����I��8E$ӷ���1��S�{�FT�b������*������xF�Rn�l�s��z�V��6}7���<E�e��h����ؤ��GP�����oe�}@���}�]zM1�!#+'W��u<GȺt6�K�<>%鹖�������y<[+|ڱ����i^����<�lcgO���f<#�o6(Ѽ:��o��̵��+�W[GɆ���2�]�1hO�}�i.��S,�a��.bXh&�a�C���wvkk���p�<�������#I�'�eU*�)�s�x<U�G�ͻ�h˭��w��s�L� ����;���
��Y�m�8V��O��������=ۯw� 4z{3/��!�/-�$�ɇFq��T߆c5�.#s��73� ��(�9�.�?� v��eH�'t���**� ��Ï��,y�c0;K�5�!s��[99��a�U�9�����ó�q����NyC�[A�%LnE�vvj�.����ScaЃsz}Â|��:r̄��Գ�Q���l)	�O+G�Fkw�����r���i4�-`�ֈ�S�uI{dh`�3r�����S�n���]�$-vbg1,���!*ُl�Y&5����)}1�[*a�S�{ka�}*{r-��Ja�J��JZ�aR�I2zY
ow����sk%�-o�lK�2���-�rO�gJa����_w��E+>����I�es�§d�\es�cl�c^؏{<��6q��	���t�i}��hΝ���ϒ gM�8�M[>{���8"0}��#�O��o�w-pq!����;��S}�8\b1,�����K'~��'��U��Ǜw6M=�JJf|͚It��q��� TY���_�l��֗Ք�6��L���'�JZ�6U�rx�=W�dO���{���at�.%�����s�Rj�S<R��3ÚZ�k~�Y����s�!6ps��A��iyhDC͙����V�ZdNg8O���99�۸����Рs�L��웍���n��b;�Z�$| �s1Pu�N��%�������F�qL�CQߩ�9��ᥟN9�|s_���c�0�85��B��2DBr����tz�!W���������O���A��ߞ����ر��������qM��s�f���6��ܔ��d�:#�ev%��D/��ku�di�~y����p��aVė�^D���� ��(�:-�R���;�2�D_
�V���6<&@����Z�Kp�gha�$�V�ő�Up�7Kv3�)�w���Bw���<��߾����v6��%�)������y�CH�6�,Gf(�O�ڷ�,�=�*L%�o5�3[;fh9��z���9��WԐv�!a���o����"8�\� +<�;ֽa�{@$U�@4�	th�-��*��v?�^;/+kԼ6\�+<k/ PK����{���ȻMd��|hF���D���[ƠT$����Z 0DVN��G,��{�v��<v~���bE�<:�k�J��P��Y4d�
����$/�L��I��QІ��K��z ¾%�w`��?>����/FB�Ӷ۫�g���n��ε�fJh���C�{���~�=W�����:@Yl�H�:��'q$p���#��N1�~�w�Gd}���zoIHX����X�ts���9Dh��at��U����կp4"�o�!�	�k�`�%j�� �[�U ⃿������1�J"!��c7��01�]�G�����Z�6���FL0��|�:�=k��?�\ i5S����Q|
p�U7�۬�D�[����J�unԦڱ�-l���v���$]��O6p�a�K���w`f����o\4��������ѻ"!M��;���0��pȧ�5�xФ���W������d�K�����J��N�<g���4i�C?pX���L@�yls���c7N�Z{��v�Ue������ѐĸ����h��-,���e�مjvQŗ��z�K���U�zv4���݁H�Xr����ӫzh�RHo)�HΨ��B��Yʤ"ׯ��TX� X<�޴�)U�^�O#��7J!��jwq���D�2���r �p���Ӷ��yq:q.�뷬0psw����n�r7�nX��b�:q�[��E.�`YI��H��:lC����O��;�8{��U���r����
��k>D���[0��'��U���~ĳ�Z���CF�yhUX��T�8wJ��|�7i�'�W��G���,�6~���춇M�m5��l�)��U�ϵ3TWW���O�L:�+�7W_H�8P�2�eH��������^i��E>ʍ�5�g�%7�CLY`��[�4�"��˳$��o��{ο��c�0I�P�����9��>� UwNE(���޸Q�4Ri4wᇞ��x�Q�W��t�������C⧩�(8h��D/��y�#/�ajy��~��Ԫ-e"��R���ް:���_���+)S����K�?z3�_:|z6p�E��{���<����0���9W�'�-�b@�� .d~u������2ܣ�I���,AM)\^U ��j2��z���2���r"�e�t�|bl�M��Ț|_���sqݘL//��ʖ��?�k�k��T�f����"��P�����O���=���Wja���Sf؊����r1��+�"��P�G����dBFK�N�8��}����G�G�ίL��,��`�5upt�J�"�J���ˣ�̵�	����� �Fp��}�gF�g���<�;�T���2���bt���{_OQ���49I���Uj[Z^�q��3��L���Y�r���z�v���Sw���K�R,p�������Lӽ�J��y���Q�#Q~ƺ��%�]N���l����77"\�&2��������e�IT�m��nz����(N��
��f(|J���C�FK�
�=?��qm���c� |@?��h���a��xn���q�V���)w�mW�E����a�X�I4��s�i����bEϭM/����iw�5#=�&��ɧ�QX��ڢ�_'�ȹ<��i*�E����&�����M(��t��]�l���m1A$����X��Eޟ�1���4<`�v8L���2�3>x��y�#l�K��x���e�3���;�Ѻ��[��Dۅ��G�B��������#�˛р~���|��4���B�<�@�jt��le1yy�4v/�D�K��x�O+��뤕O�0��[�����Zn4�۵��A�nf����d�s���(0ۮ��5�a�NKJD:Ýڱ<�=�3��T�Yel��jB��uwv~0��R'R����������Ŗ/hğV'_�[�"YZ8_Q�L=��-TWZ��F@����3.r�&�:Kq�?�{U�	��r>�7��.����?[5�V��#y�?���)�¢���r9�?b�~a�r%��Z��#羉{�s@b4әs�/{���cX�J��{��=����L��������m�Z&ʨ֋�14�yE��H�r��dvu�Ġ�D4×��`$ ����W�v�g������]�2������Q��ʉu�� �l��Tr�:o�DS�@�N.�����B��&@�ϞT�NL{����n
�� ���v.q,��q}�WV"�����v��^�¤F�ܖ4b�H�/+�]��/�.��i\�y8_8#ۑ�J�Nӵ�����9_6ݤ�290�*��8���S��F�5_��Xc�˖Cx���yoS���T��S�|�F��4L;�lIj���;��m�!"K�S/h[�=
�6��3b}#{s�o�$���Eq�g�m�z�7g�t3o��x~Q$Cղ1^�o��5���ԜOs��
�Q�:�:K�
�l�CL�-���F�4��뙹c }a��`����\���]��[ß*��������e�n;�����&3��ˢ�+�e{��xc�M�y�[�*��R�*
p�?1:�a�ů��{ʤ��� *SS	�s�hI��}p����>�NF�������vO����`{��ˏ����W�����'�'|P���G�c�^����ɏAm�$3ۃ�[h���ba���a�cq�������V�6�Ël����⨨�o(s��F5�(���`v��\`�W�(�t�#1ҷ�`���b������F��z���?MO�f����f�"ex����1~�H�˧U��)�� ;� ;��Eo��*+,�s:��!v4���2W��$:����Z2siDQtƓ׭�\V��j����vҵ+��`ڵ~�A�8>BQ�:�Q��>	���`X���Upkm4��
��r��
x+{�؏I7�C�+;�~e.�w���O���;'û��E��EBb�X!�-����}Ƚh�+���>ھ�h�HZ���n@�芜�cI	ȋ.0EP1j��Ê�����M��&��rH:�s<��3y|�
箢����˗�8\�u�r�~���q#`l`��az^J�*1� ��9H����ϣ����'�t/[�7����~��,� �l�J%o�E8��3 KŇ(�>Ɵs��ݺ��;ψ�B�����"7~=��;�U�������%���_��j��b�Ua��n*J��z����L}�k��it�y#!/����7����П$�ӫ�4��=��:+H5��8��ɫ��S�E}���]���R"џ��l��<���#}'��(:ŧҶ�f�<E���p�_�"ZB��c1��j�{�1�Ѕ�&���}�O���E�������y��o�}�)e���
̒vO��
J<L�v|�u�ϴ��\�r�����������y��1����M�!0(��`�
����K̀@:5ҲJHL�Z/���F��Gz�|��\5NtOZ��S��Q����YLP&�cP3��9�G&(oR����c�j�L�'�����S�Ç������~�;|�ȃ(x4h���"�T?��&;�R�W#!]F@�!1|�&�ՂU��Y`O� �߇���!4�>c6�c����v�v��"�+��r(���hFH�'?ܴ�%7߆�[���s�/����0XMPJu��"U�����"��<����r��"�Gwf�-�����x��)�L�e�7ۀ���=84y�1��� ]*��;O��e�0V~�Y�FL����R"Z_x�����_-ujU� ]�*EqMA�:NӋE�%h��Q��D^=^��6�F;E�!�(�]���f�X�CؑVq��6�0��]���q�P͹J�Ќ��3���1U���Sa��^��;�"�#MR�\îd��Rƕ��8/$��,���/�s͞�YZ�U �Xx�K-�oM�[�V%.�_�;���P��-��Y�g��Z���3�g��������f�.�l��������z5v���Y	��s=���%s�,P���5jf�ٙ%Y>!f5�_}/��F�>)��4���_StN-"�ڶM�B�/�>�b��Jx`4Jx�'�kɧ[o�ėva���� �wV�k���N���6�̆��辵�3}[#�7��A᜿~��;���m��q/˽|�0�W�����Zoͽ�'mՃQk����W�ڣ��H�=m*@Է�_J�/�9 ӿ�c��U�=����'�7��%"d|V�C�Ģ��{�Fd�{��C�y	dϵ�	����k�m�_�w�.x�X1�H���[-���|%l�!a]�Z�|���&pU��H��B�|����h��~�N�Y=���۶S>b#�9��]ta�u��ߌ�"���ֿ+*N�qB�RGLR4P|zb��5p쨤��ӣ�A�W`�訶�׌����`����K^0w�5�n�3�g�_(Ȟ���[ԗ+8.Z_2^<.>�ĥ�|�����^��d�94�Z�֐j!�<mȪ���d�,Z�3�Pw?�.�h/]�?�-��_+��޹9Y;�q��?m��pۗ% [¨viq�G���o#���{a{��SDuk�����J`���0{3���5����П��y��M~dd�-�m���%��Z,<���O�\�����1ӌ�
��O����!!��/}0�	�9܊,K���5�������s'�Ѩ�P�S%](E������]>=���;C���7,	,��7ձ��l��`�,\iЋ��8@���b�*�c�S�Y߱�MpXG��)z��[���A]9�N�F�|腧f7�?�9�q"��4>��g�hw'G�{���Kܪ!�Ov(o�e�~�F 5��V�D�R�dK���� <����90
�����E�)l�`o3d��boj��9�O��1���"�>\��߅��[�7�Ƣ�\�h�ԻW^�O�r��?S ����lv�\00=e\�e��`�Y�'\��D?�ITU,��Ӥv
�A��Ĭ�&m��,���b<���NLN��M��?qE��x6Ju_�Z1��Ԁ�����M@��7$�fp5�1PU�b�a	4�1�2�(���ĳ������+?��Fܒ���\�d^N~��)���_�{���ZZ5A�zM���Bf�q>���n�m���?DS�B�mW|����g�����ORRpHH��T�5��̫���%�n[���� 2�/h�����\�/1��;��+�9u-��w'�k�T�
;� C�+Y�Ŝy]�|�4vhz�@U/�ͭ0sW�-��V=(hY��x�+���X�B��V��a�9�q�?ҐT#VN��Ү��4�^���Z�4��st
.c��X,�M#�1�����g��A�w���&���ޏ���YX'}[�/�	����koj�^�<4��G����UFF�ز�}�:w/�Q�6� AK��b�~i��P�<�����g�>��7u��!a$��ൖ����i��սl�cuAe*��ٴyn�O�#j<�R��۪2g<pEFE�5��܋c�Ā�ezn,Eg�D8��AR���>.�{e�1jD�J�-����g�?�$D�i��,*�IĀat�&���+�7��;�K��bL�:�ʿ3=��'�酡��7��6l�H���w�X}P�^"��W)3ꠢ�8[}̠�p�	�g��N���n�B� +��!�ȷ��V���D�Z�M�U��`��eK`#�=iVjakDB
��>L�c?Ͳ��Z�+��1���W�cP�72(�q)"�O��;sR4�[��Vi���Y(h�8��}�+f�U��!���s�f��[K񘀥�%v�؃KF�׳���2��,K�C�C{�����d��.�j�].33CB��)ͮ??(��ׁ�-j�ms��Q�ٙzX<�	1N�1:��	{"X �:��EŊZ��
1�i�TX^޽��RH�f2�RJG��M��N|+�������!��)bּ[� �*�����lH�$����6b�`����v��,e��\��欒���"�b�Q����5�8��q^�����Y/���%2��+S6�#i����٧�QB� ��"�M�㧓�F�%o#��8M��׺}�_��.�c`̎����6;S���(���,�!�w�$F�V��h�ՑV-$��4���d��	�L��!(�ZQ��d�LҢ`���*_F��TI���OK=���O�B�YqO��+J7�>8���k��9�w��?K�G��d�
��L����H/K��Ɂy@���dh5?��}_�	r�8_�mVNU	�('E<���(?ο����~�DQ���]���!C��\Q+��d��CF��GO�7΄��Q���)rk���[`��OѩB�B~��^��q�dZ�֮ ���G��7|��!Z�!3�����G�yS2�����s�{�0C5ʤ����K�.���9�����z$�p!�t��ꇒ�1"&+ �8 ����]t_���������i)d��oB.��6���d��v�&Ϸ{6��h8P`@LfdR㎂h�O�jT~�=$
��^�"*wqm�k���5�)vΔ�#��sϢA�|�#P����Q��(0A�S��j����-d���
�����m�^x�ҩq#!�"I�	�yY1�5�0C���؊�!� ������S'u��.���ͯd��B"\T�
�%p0���<4�g'���r`P��ѐX������k�6`��[���G��!dE)�@�JK� N�S�J2����UK�U	�i9���HI~��N.��8�c@~2
�� A����(�#&�3�EB���Ք���X"�D���5����:�
��G�c�G�@?��_����(�D��J�ff�����+���8�V�&��D>ywen�u7e'?7^�EF��z�.
灓��8(9ח{�ML���KJ���m����^��]m��y��dd�Tcr�_�zU@��A��M䞿u͈�s�B�)�Uj�5�9c7:1^p,!D�_�;؊�9�)�$�|e�kw�;">"�~LQ�H���8�bG]�ک�vuS�J1�IX���km>��oK�?�؏d��S�����qf��J��� �v��cg�&�5&�tF'T��Q�}UJ�����3�ͮ��+ش.�*$pnCw�A4e���>`�?O���s�;��n��'N��f^zy��!����=<	�C�A����0=��[|�f�bε�^���~a�ʢ �}����b`Vj��,#SaI6�0��j�jDA:�5���$պ�j�H�VQ6��S�BFC�r8���%7W��t���'Ώ��7�ؼ���bs�G�#�!==��Mm==�08�����0z����:R1EW����b���������B^�俫9��zGB��������QHK�����"����(]N�A�bFV� ���R�o�����讬o��|�ϓ�d�P���O#O���6���N�^A ɬ1� ���]C���>����+*!1�w퉸��j��0K!n0���wa�&*�d���x5"��?�ɾ���� �d��%C���B�P��E�(�/́�..1�(Z��. l��� E�)Шs�(�1���W�o���Pr�j�L�ך������MUm�B��ih9S�Iq3BdIʺYԔB����8�K�"�\%(qEY�W���O1}O��s��6iQ��n!�aO�8��N�P2�]LL��Ok�l��H%�|�Q����KZآ )�!~�-L\�D��=dE >�&�
���z�4R�X;#�Hk����~�`��	n�c�'�@�ST`5���`ƾܑ����P �oxi�yj��	�7����Uw*.�8> ju`ޥIr!tt�ބ(f�>H��}@;�`�������'����$�s�� �Fñ�4��N`�T�rҖ�:HA�e����s)��i�1x�lόH<UޙÀ+�G��%�}|}�XĮ��������e�W[�T�;�;���{�:����F�N�O|Jz�u�s�L�S"-�G��o)O7� u�L��+��{	�,)��o]754]<���AȀi�n>���ΥC�ѓg:C��R�%�[�(���������.h ���ΟJ�2;��%=��K4�b6]�b��ّ�^�ۘ�S�I��0�撞n�	��w�F������5�Fz-4O��^��"O�� �U&�b����>����048M�� 9(�(V7-���'��rtd�A,�i�"��:2@O��?*�80?}4�1�OL�:р����1웾5I���o����-��9;iNނ�|����S�Q@�n��QD���Ȑ�V�����ˡ��?�Β:U�o*#��*¢�T��un%.C���!8�<��ĨSwg{�}��\�B `	��^� ����e���ތ7V#�(�����~05i�ˍ��=�D�f	gy�r�d��Wy��,'�����ܜ�����9ŷg���s�6Rz~�f�)R�4�!���<�Ӥ������U����u��ͼ�8��I$;h�e�NŎ67C��s:�6	�WY�{
��F�H�i�]�zw�D 8!����͌�֔�Z�Xgm��I���������������TΘ� ����Y�IL\<L.cMT[����^^m�M~+mo�%�x�|��R�@�������S-1���i�H;�5A��˿�%�.���	I^Q��h*��P��u���zw���P��I�!���J���)�[�����2C����C�vki>�TK�zɋ�l��Cf�����kkm��Ԭ�Lj���_�w�𫨿eQ�;��T�N����98h(�#��E�7��,4�q��T��x�0 ��>&,$�?�?�`GA-[��-S-�����-����:���]�Ht�0I�{y�S��}��'Î$�(�ѳl]�+�&�UÅ�ݾwg���d�;��|�E.2��oV��.��.Q̌�A���Q�<)�aְ�}�q!�`�QYh{���OV��<t
z���]2P�������Ol {�3��;g�E�88�����^�����Wl�r|���-9/���e[�I��`s@�/�¿i�SA���ֻp#tdR	���MZ����~m�y�r|�O#@��1��O/5��z�C��oՋG��E!ϗ��"�{��3	d=ӆ��T�%���f��䌐���7��D۔ OvŔR�.�QhC�G������)��7o݊!�œqE�O!��B��= ��U}��+z�'�^���qN��8�c���}�E�#\x�ia[`�^���s�H���/�a���~?�߈FB��O�nX�s/���=�΁0���=Tb�eb�ˢ!b��b��V�@?�_:W�
��SZon���Cc0�"Q�FW�/�����h��xN ����^}�GxgmV�����\�Q�rU q7��eQi����C�H����<)���O����W0�|��z�u}�+�X�H٢���#�L��&K��&N�G��O�}#�ɕq�Tw���T!,.gE�0p���;wnt!U��ys~����=h]\0*Z�|���ֵ��׸	���������T%�6G%8.vՏ���5��:T�Z;00P^���7:v���w^�/4Ƞ/๜�I���^��o<V�%<��mJ�������bY��Q�R\������y����� R���Y��_C�U�:�"����+��1T�:��R^?�y2��v��0��$�|�@��	^kф�-����gDB�O~�*�o�z�E����Y�7C��q&�kd�)�������O����w��8�M�uK����y/���K��{�q�쿆�^:��1�6�+��yh�A:#
��4I�����d����pl_;�":w��QZ��M+�����+Y����� B$���C,�cӽ��y��\������N:��y��W���O�.{ka�:���Ӷ��RSRUE��+��l>
A���TU9+!�O%\u�,�Qܬ�
��6)e�(����X���t��*��c���7��j��G�[�E��]�("�����(!% ��!HKKw��t� �)� "�ݍ0t0�{��y��:ι���f���Xk�g�/����T�ն�`����SB����/z�&F$z\���Rv�(H������sd
���	�߫�}qm;���0�GPf���m�ȭ���5�J��2��'��,萹�y�����x�t�k!�Ym��Q��QT�ޗc����'��J�e��-R��z�	���I>LESS�0���*zk�N�2t����h�`���*�Y59�c1[����^�`�ϑ�J�L� �/.�S��$�ZFFi�����\���}�TƁʺ�'i��l���:�N�0�V�kߍ�m�1^�!�#-b�J��S~<��7x�SP��@	i�����CD͆��yL �]yݭ�OҬ�ap��٣��9�w.�f�,<��,G6���*P�>���Ӥ��u-��A�� ����;�}+��l�a��;�Iþ��@�mn��V(���	�����^m�P���n��	:	���ݙ�P�8�{���+�/ �l1Sf��ȣ��Yg���7 �0��HH���L {��m���+O���t0����׺������5�����gRE����@�<_d�d���W{{�W䓟��!tD$l&a&y%�j6�;Bvao��a!N��Z�n��OvG�%��{�g� 
`�n�4z�1����[=��;$B��q6�t]�XR�r!��ʱ�i�4(�Rt&��>`'b��JqJ*턄�Ba.�c*��� ~�W��w�&�h�� �^^�BX�e���Ǳ�z1P>#�@�Y:����f	��G5�ȟ>���b� �Ҁ5i��~��磔�-|W��v'�>��|��T�3���ϺV*��T�(��wڜ���'�傗%g\��'l���_2�3�~#����fee���7�G:����>MV@��!��V��G��؞�c���lo<�:�L.(E����{ hKƳ	�ד� �����X.#4Ǆ��ɾhB��v,^��4%�M�*G��Rt[fU�S8���	��Dl9��N҆������4����o�JW�a��	�� ��$�+���a���^5%B�Z���0�)?b��D!q�<�Q8 d�8����Qզq�å��k�"7��7�#PʫU���5A���[+S�����gr���T��z��Un�L+��������X0Y(A�QS���*��<qֽ��)����Z��jA��hn�d+���hQ�^^���f+�'}�����  �� ����np�e֕b�8�A"&����BA�L�o����'_0y��ԧ2���wlީ��i��Ww�\��\��}u$�"J�w�'ӽ|�x�O~�=�Ŀ~�w��������Kϕ�г@��\/n��;�}e�p���#a4!\�3�T<yB���B�/&b��}$��#Yi�����J~�M�G�``�dE�+�O�e{Ib���<x���O#��E�OH�F���'� �v����u'���SEE��؟�ᨾ��(#�Gӟ��r���zv&�\�{ E����1F2�"��'�:�TUp=f����H.7�݉�hL��y��Z=��DOF*7yΏ���~m���D;L�͢�$#���q.Q<u8�qɕ_�a�M�N��}&wi��:~/?;�`�C�fӢ��V�ג؀��ф�7�
����ި�!~���QO��0����Ȕ���ܻUf�R��)u�)��q��s0�z������HK���`I*P�M���8(�����ex������?,`��1_��g2��oͱ��}%-�~F��
� �1<f}�7OȤ�����
F$l��$2Ў-��N#A�Y��K������A�9�w����v�g�Z?]�\/X��7�QJ{!�h�oP��E��~Rc�uY|�d�h�.yh��(⽓g�+T�>Bt�0���;V�����#���b�����)b�C!CHҤz�����w�a��m����cn�ݷ)b&�'�]}f$c�?�f�<�N����(�
Ț�!$Tx��-m�k?UǞ����]��~-o6o���(ZBb_Ǻ'�Ѭz>h�k�(����˝����f�Mz	���|II�S�t��%{����N��nBy^ �ֺ�)/@�3�.̯x�"m��;a��r�(�#^� #i�wN�M?`�w'�;��l��(��>	@�b�2�xg���zx��bR��+�������t$ �V�#tDO@�3�w>6�M�kP�n`4�����ƣ	E_��;�o������)H������
�O���t�;p�J�I���^����.�|C�8()�翝�B�J���6-j���L�O�u���Y�N�%Lml�x4��8�Y<���M����IJ�l/b|���4�rTLeK�
�Q3�LU�A'_�� +9{�SC�Q3S��R3��3����1���3��� �>��y���F�+�ߩ��m�'+�� )��oC?�o2�P�t��٨�v��{��*�wh}�����uh;ߠ?�K��z+Ѹ�_@t�HH'������;C��h�G��_r��A�@��Ē�"__����-��f"�!�2'&�fZ��|���7�y��������X)c7h� ���u9�U�|�~<X L�����5X=m�n�K�_O��_]wlS��ym�%�rzdu����ߧŨ��g�4�A_r<~�?��F��"��#�௟�y���l��y�����i��������[�h2/^�#X9]��O��x��٠��봡u��ww_� 	+UL[�E7A@|��nI�nPd�8�k��3Dk��f	�=~�-(�36=A�_�_��:�m�\�m5�2=.��d������.|�r���(	(oT��&�^��D������iK�ϝ.����r΍i�v����`0x��B�|��Zdu�T�/$$$���QF^�:�]�V���%dݭ�YBqP�o�5t��M���΀#�w���xM�Ƞ����ޗ)QZ~�T$O՗jY�Y?E�WW?.~�7Iy)�<t�($��~�5�d���×
V�4�F��O��?��ttԻҝN7��B"��r�s���h�d���{��L=S�_��T�|�E`��+����$�j��D�ꋦ�\�R�]}_&ItPS���HT�8��ؔ���y9>���9[��33��~	�{�B����Ú�_o�o��G+��p��t8ҝr�خ��w��{����+��-�?͝RGL'�wO~eh�Z���R�Y�.�`�� <G�}o��p.�]�k���bM��y	y��o����(C5�����! �(B`зۇk�W���dlF�p�( ��v����{��===YkkF���4h
.绲�./�����
��xo��CDa��^����b�(.q\��O�������-<z��vV��\ߢ��G����PU�~��3nP�`�
	����v/|���>x)��|Q؊������/6{�wҞ�Gr����S^�J�����˶Cmly]}�Y�h"�������&`��_耫͂c���N�nN���oJ�0��,�{6CS�	yw��^��?շ�����eZ_<UO�-���+�-~ƿk�'T焘�|U��γ������_�n2�P�^�]�g0����''W `�z�x9(t������Au����3L	���3��
y�����*z���b�����������S#�ov���^#1���z������:�o�<�ݧ^o�����*��ZIb��%�6�Ҭ[#��55e�>}��ȋ�/X	��@��S�5bQȒ�JI�L59�$.i-s�222hH�uZ�í�E�<=j��)o^ņ2E���֋�޺Z���0c� $[h��v;G�n܇Y�jD��I��������H�S t�A}n����)�KcϷ���H����k���Z��7�=.�}9s�H}4�)-%�������׹�f��Wn�tOw6����/*y�����a��ޜ�X V�a=b��ۉX�]�,2����O���]��srp��:m�[uhI�62�������SR�>�s��5p����bRIM��^�8Ђ�ۛ���]`���hQ777�����6�̖~�"�5@K=y���_�:���8(d2z뺹�8A'�0��u�֟�A`��&���D|�l*:L:��k�?�������~kpB���[ǹX�F������R�iB>��)oZo��;f��u�Q���Ʀ��!��{��P�J��&"oն^�$v���o��?&���J��2[=�����8tp	"-w����tY���^�����b���������ȏ��������ف����-�R+�.��h=N��cP/J�qx��ٹpx�r���=�JR���=]������ ��낒�.x�c_ �0���*�\��4�;��MؓsJ�`�۫�[Y��/[�N��ۦ�v��󟃿��̶Fr�#)��7����xy!�O�]��yj���y��ˋMSk�Jm�5�`�^"���P�m@}��ޛ���l&�q��h4����s���|���CL�}�` �{�{HOW������.[���.ބߜն'��{�K���%�}:������N;GF���:�H�u}6k���{���֎�.�SB-x�zt�sط�P��o���%�,t�Fs����|�3�d��l��ϥ�����v��&�����ԣ3��M	��~��^��n�䓉j�c�'�>�k�js���:߄˭�uz%�4NG����$��z|"�B�L!����:�A�ykg�������ь[�)�7��t���ƴ�Zي�( �K��8,Z̽5Z�^F��ʸ��n�I�:?t��9��l
S�I�Iw;�n���u=Ȝ���v�Nؚ���<=G\)ؼ؛��׆
��"����Қ���.
���!�O<�v/m\��jMN�z�oW�?baa9F4

�`�4_����rZ��S������.}�(��,k���}�*��R�����d+��Q멵i�g'S:��4������b"�M8�����9�(����/�P�&�>!w�B���8m�a|9BA�����}"�h���"R��=O���)�Ǆ��+At�J.�������@l��7��U�ʤ����>���-P1�#�iP�����k�����5M�'�J�j/?�l�ϭ� �&f�Q��.+W!�ܨcI\L�b;d!�̧���z�����a�O����hF��ZO�2�f-GɘS���Ex��%�s	I<�"�o��<��z�o󫼢*k��
-�U�9D _Bz��h([��>V��1�g�u�G*;���)���8R=`�߯&[oT-k7����8�A�p[���V�s�'�f;ilw�E$�o��S��6����5~���\�}�����zad�?�����U�x��WED�y�M�r���u�O}nTR;Ӏ0�i9%��R.�:	Z�ɪ�^�4��Ӳ_ձ���ī�k!7X��{���$�=���tc�
��Y:��u��g��tY(�kw#��C����B��5���G�Y�,!S*4��ծ����&�M�֫�I���S(�5�I~�w����X|;���U�$��)�l8Kbtl��Q��5L7���S���J���\_S���{��7kkv�d��M���?|��^Y���N�"�T����>eD��3��d�1�3H���u����n��V���E�Se>�PT��'�&�$�˒+%a�Z�ާ^&&&��n��/�]���LY|{]�~��!~,2�!�)�9�d�r0�d���j14�"��T���w�f�Eg���@�[EQ@��N���e5ш�徙�R��$@IW6�lq��}���2��H����ل���h6%�k�Tg>N�
!Y��m%��hk���I�r�5��ԓ�=[�Ϫ�0BNʰs	�>��MK��\�l�b~xʔ���"$`2b��g������eb�=P��z���A��Q8|�����W[�$����ĺOK��$�ރ����@���įK������!}v>9������{fC�"/�.�ަ�v��t�R-T��L�{b����X��j9܂6��`����'o
e��o>e��[x�}���ʲ�P�B�?ү�h�[���Э�e
��c�Ľ&N��i)����ZoK)��g^���*�n�C�2��ڢ��{�6��ZO��H�_��ʫp��"��u cZ��%'ĶV�@��*�V�\����b��FW��o����̒|#5�:��ǫ]��b����o_	��e`W1����t��N�C@�%��#uŹ6�b=�|�ra��*��x�����	�6|�;T��N���b��?���3+ �Pޯ�۵�	��������Y�%/��r���������v��1,w�	cI1$vE�?�#D�<~�35��E;M�Y[�T 4���u�.�+��U�+���MQQ5f)b6[u����8-�;hk����r�ĸAC'�m#��)�o}���O�� 9��Ƽ��)�t	 ��4��16�4��N����:k�{�*�:��Ǥ6�BB��\$j2��/@G�K�F[F���$�
�-�$T����̛�X�~A�k���7�qmnm��m��ʰ�	�9ۋTD/���Zof��e�O ��r^�P�K������eb��_�J�S��A
��f� m������3�}����o���[:bl�e��ҥ��cݳY��t��oG��oA�������j��ZNxUe�x0n�n�/�Y�M��� Țo�k�'Nv>�lD��}�M�x���|'�n�5i��@������KL�o~B��u�������˺��P̝��]�T���ٹ�4��a�޽{S����s��ò��=�E5cN��3��V�d.����͢]�7�F#���E�}zP�c]��Wg��U����G��/��c�4:3v^�'�`?-��]���l�ֲ�=|��U��6�{Ȓ��N!=�{�ZЎ�Ǐ�2?�l��b� 	EhT� E�l��~ aymH.\��YH����"��K� �G*�z�E/F
�|���� �bb�q�l���BU0�t_�F�;���8-\�P�K��%�|:?OOoNlډa�4�o\&�hݤQ"�����@N�F��8��a�*l�E��d�O�d�B"!N�w�馃�� ������
*��;*�d�m��؍$�h��n����$%J��=��J�m(Rr!q	������xS��L��k_��k�J\����;�s�>�}�O�I��ݟo���Fj����~s��k��Te��Pe�; �jv-��]I1����V�n5��O]p;M���Ej%ݵ�T���Q, C�Zu��nt�Q�|[�<MZ���]�n�u�Ah������ � ��+��$i�zv\Lv|�J�HK�*���Ƴntm	�LZ�>���P�n]�j�l�u����S�.H�ҟ+Wp�~�3U�j~�����-�������r?�6�i���4������zB�'�y$�ګg2���c�v�b�����yer���`���e�A#��E=($�  bV���f�f<0���ͭi�>�b���~U�,f����T{є{�� ��������XB���C�Bڣ'�Ņ���Ƽ���*���pG0���:*S�Q9��MU����@�B����;b�X?ArQ��))|��nhRYř��+��Dz!j�t���,�[L�]�����祱�}�[�d4�ݸ螚.\�?��� ���,��X�&{'����=���@�P�n^��#�q�����j���S8�4�vmZ.^v�J!����0������d}qk4OQ�S�b��r���zy��g��%Em�W������}�8�	<��u{���S`�n�T���v ����FB�ru�f��!�Z���rEK5U���w��kڗB"$�w���	V#�r���D�:��q�1a��������b�|�ĉww�W��l��C�.l3�F�a�>�#��B�Q?�|�+NƤ]�y_����T �/���*˸7~Y�b��f�A�I�l���}z�1����a˨�r�G�4,&�Կ�#.��8��ĹE�X��p1kOs/��Hv]���a�i�3�r�1G���͟�/�b`�Ѝ�靜+W�b�,�`��?��T]XRf5}Il�1^}=n�mȨX_f#�`l&}D�5��Dp���_���� � �ّ�����io��haU ����P/Ն�c�'�.�Q_'	xp���iW�dK�:���ޛ�r�ϤY����-|V�_�s{����t�������:1����8̨�݀�苌�i�F�n�@��S�8��	*�O3�û��F4��̕'�>g��߉�,�����^�[���+7�� |Pk��ʽ��ݶ�5,��X<�;�ɍ�t
�����Ȋt���y�}��8/��J�W�;�s]�g�)��/���Rg�v��Y�K�ZK/�"�M�����u��KK<�Y`>f5	�Rమ^EGؽ8Tl��+v�4 e,9]���f3�u���fc�`��A/M�H2>�f�S����f#vr^Ǯ*�k۾��no*"�W�4mxϤ���Zr2�%D��9��2�$2��>_QQm�;���r��㛩'��1q��oY犟�X���˛@#I8��\Z���
Z�+PF��0�t�ي�D�Wޓߙo$|�i��^�X��+�Y�d��Օ>|��fѺA��4��w�3s�m��F��eO�ط|w㤘6uuu%����L�z{cϛ�Mz��}�_k��3JGS�?�&㴚ɷ�8�ɒx��o>kĵe�C�m?�e��Q�0�c�s7�^�3�D� �����R�OZ:6 �Vu�mzQ��eD��9Oc�{뙸�r��������n����^Q�l�:���.a[G*6`��Al���W,Ѿ����_�������z5��D_��x'��H�i9�IRv��y5�@'��o���p	�0�}n�	B��db��3H��J5�5:�����R^|�Ӛ�4g48V"�</H&�)| ��p$[:�0�C��"��*z��|��&�d�aC��=	�k�����{\Rr� g��E��Y@R*d���*U4�mP'd�L�	U�t�u��oU�vw���G��j�{k�2�aX[[�]PsO�2	;�
v�Zm�fZY
k�8S!�WY�YcY��Q�b��!��ϓ��.O�GW�0���^f�o�_��=o���z��[i1Y�����ݸ�i]��f�>��V%�k�t'��"Dd�e:JԾ[&�EOK�tk��vYtt����JY���6�w�^(�B�k�1���	9�(���5��&�������\m�����d	
�H \M~�Q�B<�(&� �1A����� ���+��/��ۍ�+_ƈ<L@6,�I�dpn��Ed?�(#�T��dXRm�F9G��I������f�~B�H�?~�7�o�8K~��V���&)t6�����t��}��]W�Ը��-#)��(�5��,BcX��V N�w ���@�a)\6?�~� �LO�;Ϗ�����h�6.,P��&�	
,��D?�����rø�F]��h`��Ɉ$����pEH��c=�
i�"��||E-�@xuL�nɮ��tG� >�6�8k����Y�t_�W_F����U�/)w}i:�nQV������5))4����5x4�l�L[�ɶ�(�aұw;z,F��@L0���R ��;�s���N��;*w������*�?�$���ӡ8��}�Pe�`�oRR��j�os팷l�J��DX zm`�v�����~�yٲ��T�T6~36�i���D|ZH7Z��� �@PQS|�@>��*ƶ���"92ä� ��mS��$����^RJ�/Y�^�M����e�;��h`����Q��������� @�[�,P�+�.�B���}c�Bp�[ÓrmrS�h�R]�ɞ�n
7=����$6 ����%(x3<M������'�����5*������Fw৹\sO�콼wѨ�N���%�oCD"[��|M�sÿ���)����AP�O�]]]�[xF�{EPF�W�!?�/M�n��K<U�#,�=f7S.�f��J�]�ea�~�]hp*�w0�W��H�҂mh��?�6��� ��q|��ԉ�Y�;ã��L� (Fѡ��_k4{�b*TA��t�-��PC/����K�v'�
���+��R��懁,L��N(	�5�]95��H�,!Sm��u�8ƍT5�J���������#G���9�Qd��M�m�A*b�N\�<�he�j,ݴkj��?a֓"���*Tt���g����‐a�?h��'���H3��a�e�Of� !CW�]����[缛L�GE,�\*M����Z!���g�.1�M�!W>^����	I���H�xT���Ϳ�j���t�x)p�'$/�Dᜭl���"��Gtn9;1j4�ό��3]3W�
��7g��+���8�]�u"����Y�1ۭ�ǡR��Ŧ{���쵴R��)�/E�|�����܎��^�ݣ[<���"�?3�� ���{�-����
`+�.�h���B�򮖼q��5�я�7�./�������/�ܟ�W\/Xi��G���h�Y�O�xEVb�Q
���u/%t�m}���j�z����ϵ��s;�Ƿ�W!�wu$!E�No�A ����;��f��c��޹��4��X�1r�\�/U���|�=���n߻ɓ�����KѨV��/7u�SI�}���>�c���3t�<�*��Z����Fk!�A����d�G!����h��[�{u��p��5�2�Q���@�y��2)�����8�(��Xd_&-g�D��44}l���0�xm9_=�"H���T��u�����A�]�,�o��p:;�O��o[w���ivx�e��K��XAA��ϫ���Uf<G�ud�v�n�^���7.+/��i;�EѪZ�<��=Q�۟�"���/�v.�xO2YB�tPi4.ӧSA�)��QW�iqy?�}A���YB���m���c�X��uֿF�%�@���g���-X]U����8z	G����M�o�-w��l\�70�R��7^�-`���jkk�>��]��eNVFRO��6�
��L8�S�i�K�s�wF��J��x�@����ƣ�<����Br"�q'��4��P?���y�Xg�����V�aD`Ќ��QX7����?��+�x*L�J���� ��/��&�;��Na��g�&'�'�h������`r͛?�w� Yc�{5j�0Xs/�Գ���8b��_W?�չ�F�R6��g<�c�s�.kj�M����s��m�Q�����Oөe�湤-e�z���>�����?�G�a��!��1���x7�x����k��=Ryh���CpI"��^�J3ʇ� ���,�����?~w�T��WC:�5�]�����~��5�LP}�X�q������A��}��C��?�`+�p4~�}�^�Bx�e^tr�yx�.�m4{𞏜�oL��k(�:���Ma��Q���TΒZ��j6s�&K)8Gr�rO��j����A?e����?��{Ɗ��l��[���2�����{�}�ѩ��y_�Ζ�\8Ygо�� > �f3};�Fȴ�$�d�j5���\�4ı%���l~��$��g���������
ꋶG4]yT
NkT�C=[�xL���b,�Fa�/�������\��/��1����x;�s��+�ne��}ϛ��ڣ.8a��������˕�8_J��\��Bj^!�Y���7���uO�e�!-k��Y��?�7��?�͑G΂��P��ݩ����d	ϛ[��.)=a�k̕iPB��$��~�|� ~�����j���K���(�:#�cj^���W)Wc���=��3� C������s;l�iZ/4������?_������0q"��4���:�cn�ڕ��/�A�?�������#)f��M���U��0��c�����c�;�i���"�YP, C���6�7�j&�A}�~�ǽ0�9��ڏ�r��li���sԡ���/-G�¡c+�X|0g,hn9ɹ����4���y�T,㞫���f�k�����$���C�ֻ@��}��r7��1d|WTTq�{���#6��,�C^����TJ�� ���,%o�:�^��/<&�]�	�	�����<�k
��~���"�7XL�BY~ �;h̚����g��I<M�^_�S;��-�����a:�0��!�js�� ����b:�z�n�B��ץ�*����@*�T
'#ϔP���ܥِ7M�l1���d�;!�@o/áaZKY�x"�t-W��}�����83f�!KPM�x����z�����+O~vw���`��a�v��(I uB@E#��W琝��q��7 Qʑy:U�(��&��ş!^'��9�nLq�O�G�-��vL0��t�ԇ�������y�c����s�3n��Ҁ�9t�E`2�:Ѻ/Y��X�n&u��m�Cg�R�L��B[J�Wt��_@
�_��K�}b�L��9311%�:������	��)l+�������3KVm�H���6�<?+�$\�7��Z�0���bF6]D�M�Vw�KF�%�I���z����R�X�
E�#_.oX�m�s)^2�������S��̞��l�>r�W�@މ^�h����%O%�cq��1߻bw��v�g���O1U]�H�´�Hy���6�&JuSȸR���:z�k@�:�2q��\^���u�h���o�o����0��$�/�jm;M���ѥ��OV�����R�$KUd������k��\9�o//�"8����H�
��lS�N��x�V�����p�\N_�q�K'��c8��7 �Ę�I�K�����-����ka��ƺ�7�cq��[H�(E���Tnz����՚�]��yʬ�?P۟�'�3���A�d):��3F��j�O��+tN�����_�:yM���,�##`p�R!�fe�`��"����"��e�j=< k���ۗ�)��FA]�(R�j����-ܬe�u�m�vR�����6��$�u٢STlP������L��t�K�Gn��5yrL���O�2�P3���N_����Y�G�3��y��=�l��&J��׹g�-�ۼ����KH�����5�ػ��ɨC	<�פ��� �zڕ�X%�tV,�z�e�3�18��!�1z�cc�s�RdX�YЊh�	���2����A�$�VH�Kq�^m�>�j�o<ŬS��r��F�Ͼ�����Q/U�C�.�!� Tp3�Va������
ɸ��v�[t�Ekmy(�bZ�kڊDH���q�kZT�W�g]�yb�r}J�u�s_yos!eD�B���>#���b0Z/j����.�n��j��k?���C�-�`/�߿����85u�+�ӫ�~�I�F1����[Ed�g��\��6M��Z������rtJ��'���MQ�J�#��'$懼�p��xM�5��)�eˀq�G����i\��<�t&��]�ۮ'l}ɞ��������~��<����*��X*t(�|��Ko�=�;S�Ƌ�![5 �Jn<�[�,Iy^�E<����3��F����]\���=��f�c�M�x����V̈́�w�@�S��M��DVx?��<V��$9�d���H|����~���u:g^�Gv�L�)i	����w;�!������3��,y��p�s�Ỳxlr�g�P��O}i|���D�\8�gTI�lon���$��%W�K��ӛ'�"&m��]��Bf�G.����r"EK��v�{:�W�1l	f+�;�+��ߖP���=cb�~�5�Xz���]�.g[�c�
�6�W�1.^C'�� �v�f78 y�������f�#8��R�����=�p���{U�4{@�B�����"�F��'�����h���#s����_��ymb�$\�&Y��R�ֈ/��%���z��w�$�P���P{!y�O���!z���&}J�3�O�{{u.���&>_�9���]Z�p	 w����W�0%�����H�B�h0.�9�d��|�T+��iS3�b��
j�el;*��ʏ�����H�^N�Ű�vS��<@{�	
N��L���zp�)�ӗ��cI��!wsXMYi\�k��y��	C�NH���,�:����"k���g��5}`�q�����Ma?D�R��.�;TgQw��ܦ7�z��~mrqٲ֫^���q�m!�&�[Ҫ�zt�=E]���D�P����o ��N%`�
�]_�<�oSx�A��:+bL��1<(��F�}���Pn�L���!����t���%�\�zyR߼����T3��>l�BU����wl��nT��5���Fٽ��2��5��2�	2<�Ĥ拾�x�����.�F��n�H�����Ǭ��b.�zv�ߞJ��蜕hV��zx��Jg�`ʑe��S�l�hwd2�˨��	����k{N#4a_Ⱦ�����%���RK����q����6�}�	��Ǻ���g�ac�R�}D�Tm���Uԯ�_�	}7�T0�I�g��.vڣ*�!������&��j�>a5���A�QO�e��⃙ӻ��ְ��Z���{�ӈ���I��_�!�Èd�S���æ�_LZ����.����zx?��ɑq�&�l3�B��9hj̆&���}�dD��h.��KDj�K������p�U�]P�,zˤ��{��f빺c!��fF�#�F��N����Ǐ~��%)e�8-bB�Q�����8Qi�g��i٦��J��.�� y#���������y*���G�/@J�3E"y��Q��j��G@�J4�a:O8G
��^�JL�	����&}�7��Ґ�	�tL�= 0�^�����L�)� ��k]�:)@N�q��zR����P�b�����:+���t!�����ܥ���W{��R��E?#���x2q|!�2�+�s��l�/��jge��r1�j���<_��Z)+=�Q0v��G&{��2D���y��EL��(��o���́T��s�F�]�y2E�[p{�ݱI�F:��Τ��D�����"ι�:^�A�5�GuD~A]1]���kl��dm����I�r6{\��ْ	7�.���l�ӢdT�|0Z���z;}U�Z���z���|�c�薽��͇�Lb��)�<��>M{n��$�F�cmf�]{}�'j�h%x��ȉK]q�.��Gwr���!�ƨ�C��O�o�Y�2��hG?�ؙ���/._@�qI<n�;����4Q��I༅���$ƥ��>GM[nu_�������쑦��{\c9�F�]�L�`�m\���8(�J�⣅��S�Ksw2s�"k�^1
���?�Y!�1��'�λ!��B�o>˓O1!�1 �X�
`�BW�q���7qKRE�Cӕ!��w��Q��`L~��w�,�ݰ;�ȉ�Bb���p>z@�ލ�L����z3H2�_�^�m�!v�2�b�����˼F�K�}b��u޼�BGĤ����d�K9FPW�!��:*)��{����˄�O��_&xxr���a,~%)MQ/u#RxLd���S8����Lƣ��QL�H�2�Z6`����fot��-mk����`��T��wJ5Ftٲ)�=�J�`��/+gi|h�����~����8�a��B�n�'���/	�$���<.����}������1�����3�7�A]gT���U�ᑚU�ѿl��@�a_�:�[|�qp�z�ܣü=g/vO6���0��$��T���p�����6�\�;L���= S��mx�zY�J�s��w'ݧ�'&�|Ƭ�4�f��mc"߭ǅqZ-跆��	�Į�?��իF���.�m��f��̐�k�T�g�����pP����Vm@���oiC���@s׾�HB��&��Eeޖgw��QPWM�E&U����tE�@n��-��|���7���.�iT�?t�A�Sh6�M�r8n��%]������hݏ�:�+��|Ʋ�)�}Vk���]�P�0g7(���a�����4ˌ:͸

���:�c���4�lx*�r�3�_��{�-�O��R �p�&n�0�ӫ��;T��[i�#u�8�N�)��Ry��.J�j;���<&��N��+	�}֢�`;FH�B�Keھ^��_uAq�1��2E���B�>�L?���q�`,A����Q���K�M׊�׋�Us��<�'���,��mnXR�S*NR�.���)���n�V�u��`!_�B3>n��^��D�/'��'�D�����E���`d��mġ�Hh�˵ݲ2m�vs��`P�����YRoGݎ��V$`^����G�z��Q�ѓٛa�f!�T�<���^WΣn��Ԣe�ͯ]> B4�"�߹7{�W�[�_����fA12W+��p���u��8|��e��f�H��A9?��;P)�M��N���U��@8v_��D�����X��ބ�f+(�@@>�*@�	a�ȱA?������Iy��{~T�V�RC�Jci k#��h ��}u�_�:H�c �r1��LV��\������v;��=�V$R��B�-H(������.���X�b��ؗD�s����$�� Φ=cg��<9N�&��]��b���4�6���i��<ۡ��wj5��ۓ���E�m���3�(�,[֖B�H�Ъ���A�����Fc���S����F3�Kf�G�����~�:�:��Il�r���F�R��F�����軂��Ϫ3���tl�?{��
�"1E)ɧ[�`>�2f��<�S�MYE��.����U;z\O�$��&Q���#�����k�`��l{L�B���p�y��X�:��Q�Ө��C[�tt�[�ڝ�H�s���d���Q��6t���}��P'�4(������g�X�d+�&�4�	[T�t���e|�j&�4o����`͈1����g���{W�3�wk�ڙ�4�F�+�"KP}Ju�C�=�v���Gf%��O��^JU����~�����*&s�>����-�YaU�>���ϓ$��ް���8�yp��T�M�o��+u�s�F{�\A���(r̮�Uo���/`"J)�H��)��tw+�H,-!�% !�H�R��  !�4,K.,�[��<������s�ܹ���ܙ��|�BxN	�,�.�D��h��9f�����Y���V-��M='�x�V~D[�#��˗��l�P_�,睤�i�k��c�ۯ�k�	PP���+��ގ'*�`vdk�:��=��X\f�E	�����Z8y�p���z�.]�H۹nI�KiD�3���ݞ�/��`�T�
L�ufa���!��p�!���k/
�����#����5V\�{�5���v�u��2�o�+��U�~��ܼ]��e��c�'k7lUN��8<|���k���'6]��!b����ڽ��L���ޞ�'�\sE|Q�P��!,p����i��j�%0f	]���	VmU�m����f_�M���Z| �9�A�:W1'���8��_��z#�u������/����Ɏ�|��9��ü_Z�}������cf���, ��V�X�Rz�[��2�������91�Ma��KS���A��iܒ8';S�����v�n��u:�x��S��Y��!�]���E�3{���u}�h�\%/�TЄٔ�({���+�Z�/�����)���*�^�9~O���}��T�f�q�ԕ.�U1쵼�-D]��m��̲�<o�i4�N��㈎�=�>�Ż�b��7g�2OO����4�g{c�̙ܞ�Z���~��ow�Z�F�8�v5K���-g�Ѓ�f��b�v����s$Ni������í��ǋ����ƻ��}��$�1Ii���>�����<�Kռ_�(r�BP��Q�)�4e��HHֲܶ]���'1�<���x<�����>�ƹO�M��"6M���ù�~=:m�bC�����FK����g����x��˚�gwsz>��-ֈ����E*�Qm���7}�ġ�
5���ih�4���㛘��#�`�\%�
~�����[2]a�!њ� ;ϗ����������o��0؏��U�I[WH;�/aL�8��E��@�F۝��V��9�V�����JG�৭�����������S�� V����=41�xR�b���M�B�n�".�K[ˠZx�v��P��x�%G�.�35�{�噮� �?����Vt������6�N�3��d��y��ܪ��B�?4����&q��K�7�o)���������b��b�����Yu�����hp("0߀����|����JXHip�O�ݓĨ����g����������f��љ����~r�f��f���=hZ�)Ү7sN�8�!T)ȯOe㉃�'p	�����W2pҌ�%\��,۱�ޛ�b��r�Y�]��s�Ӧ�"L�x��^�Z�,�0�;��?��/���;��Ȣq�T���?B��k�"zW�())ݑ��h���k��O�����K46�D�n�u ci��,�^	������y��
m�'��6�~�����t%ŰȦSK���7�&*J^o��6w�9Z9��|�`�i��a�S��3�"�g@�L�p`�vA�`�Zo4�3�C�'�l�.��cG�����Ic�]k����ₖ���V����R����X��o>�q��7U?�	Ɨ���x:W�`~�ПC��Q�5��Y�~�e7wgtkY�+�d�۲ל�"S��?Oy)v��6���cǚ5b4��g�z2I�0[XX�	Z�.�s�h�jf��Uq�Y�f+�h�;l5��2�-�������<�˕$5Ln'@���Iу��6�ɶ�zg����]��i����?6;��M��1j��6t
e�����R��%�{e�@_�:��	���FמI+�'ea�U��o^`��=|*u���aC`�l���<�Ǚ*aʪ������$������e�i�YF���n����Ӏ	��a�-�˶���9���K�M�PZĲdҙ%�v=�)nd���/����ӣ�E)S�ۭ��d�����.W��B����T9`s���4t��V"DLޛ�Tݎ��_�±=7�
���~:�=W�N/Gru2�T�]I�C�V�	�5� e�%�R�0��<��O�'j����w�>����Q�?�n���ȭ�x����~
������kԹ����ƏO,V���
�f�L�Î_�!\]>�6؇ۓFi-�$W��t����Т�q����0�C��s|�>*�-)�*��ŵ@��E!�NN�\`_�a7�(V4���SP8����c�f�x��JڣCl�x[e���>��"h��{�[����r��\����\��M�7�"�tX��`)�!��{>]"x�_�틡f�Ę���+��UE)=�&�]�V�v������ek��S�3��J��x���̮���!�ڸԃT�g,� �#��b�Qų�gQZ���M�--1��:�T�룙F�^(t����l���_�_4��d���r0��m1F,�AA]HG�~�)Ov�̠Y�n4]�y�n��ZO�����C����Zn1v���8���[�;{�u�=��N'��܎�j�|�|���s�W	a�(ԡ�\��gyU�(t�!���u�j_"�4���k��=�8�WH�0�x�c�0�7�{�q(�y���~n~�~��r,�v�T��h[g=V hMڪ�w�(���3m�%SL��"y�Wk�)�n�X�'�ЇI�y#Ah���E��n���ʔV�̡��A=�%k��x-sJN�@kd[�?W�M�j�!��&��^?�xR'oN�kJֆ%N-�����c�ki]�(������V���.�h�}��ZM0Ud
���	���+/�ޠ8�EQ�������e�[<��6"�DȖ}P����I��b˹*z6�ԟ`�X�
m3B�A#�{�����*����n�i���v�w���p���i�2@�<�[Y�e�b��T!��=�˪���x���7���5��f!���#K�Uռ�<ݑ#��4b�"�ebxB�=cҡ�E����r��|�q�q�$�-*Q��_
\�8Ja��E�s�F-l]8���;����YO��M�z��_|ml�aw�����rw}zi>wm���i'*�.�
�*^24���p�.nUʥ��O��.r��G�&��n(���`DC�����L�_�h���o��:�>�)�	�WH�1j���:�ڙb�6Y���&�*�������t֕���m���� �
J��z���~�8l��m��>�$k6X4��L쁙,	GT�����.�7��6���!~�yH�m�8ƂF��d�?Rh���|�2/jf�Ŧ�z!���䲫\a(>����)���n�Th��_k9��h(����c� �JQܫ%�Ѐ�o��#�y��&�%e��������PZ�0�7񷪮��2`���ݤW�zp�~S?Ԡϲ�@�J��r6 �e!�^���sQ�w��C_�/oBH"k��n�G�}D<�Š	�xIQ��:{�rpb�=O��h($V�7�v��ٵxyP�d�*���q��m@Ge�L�����MU������[<���)�¹�N���*��&� ���d_�ߥ�)2L��8�Ԁ�>^�+t7��rD�����k?���0��p:u����>V��y�,7Gҭ��Dt ��}�8<ƇW�k�{VI��L��w��I��C��۞�]��P��f.�,�*�9���Cu@~ ���G'3��*O���7M�yeYx�����_#�I=�(�M�BN�M��R&g�%M��U�z����Q۝���瞙o�nN-Mh?JJ�wr�銢V/j@;Ѣ�C(�\�gS�z
��nnn\I��E��}>���Q�se��#~���nÅ�tG����������*���Jh�LL+�5zL��	 �o��/�-_K�_=��M�W���sQ0�4u�Gz<�(?�Y-�����H�-�@�K��D�#1�X�)b�f�[���/F�F��m�\���]{k̒�"��C���{d������;
��ϥQ��I���ޓ�A����d.~������}=��kG.����Ơ=����UQ�r�As=��O���|�S�yV�:])J�)�+�vSN4�OK��{���@#N�Ufx�"G�+��3�av�����"(�|
�������kTk�z�j^+��%��!hx�A�Կv�5 z�y�CB�w���
ݪy��;u�j���|���X�l:��o*��.;��e��DWB(���:��X���c�)c�X,[|k��z����,'�.g%�OӬ�R��Hs��$߅t�+|W���F�gIܛ_�k�NU�2�Jl���3�d�*��xl6��@,G��-;7�5�9�h�G����h�jNE����V���!]Ap��#j��R����)_�F^ty���z!~--�G8�؍��Y��ђ�8�dv�O�����`�+ȫ16Ů��s������7���A�z��I5,"��Q1ˤ7*�=�^����:�/d�
M]�J]3ez\^ȏ�{��ż63���Q���+�%�5A��w�'���!?��O �R��o��w"w�]�Sc&;�β!i͞�r[XD\9��n��9��am! ��	�뿗Է9�A����c�#�X��n�0R1F��Šѥ^7�j�*��[��J����Q��K���A�)z��I�bxt1lq����ݑOρ�V������x�d���$A6:b�G'm&Х������b�����#gQ�Mv���b6��mX���F�?$�q�9V�ĿiQ���j��YR&2��&��+3#Yx.L�N�A��P��X#�k>*2��aBN�)�qIj�H��QaTI')��FOL�-�����D���7q_T��V��1�J���U��ꯛ���K�^����櫟Jgo|����I8 K9��_�T�2�y�f�Yi�������E-�?̋z��S��{09�Ė�AAjT���A����ܯ5N������;..�?�fK+"[��#�r(�n���L��Y-A!5��#���(�M+�@��ޖŊ�8��7p]�jn��_fKE�r�ɣ�OP���nz�X���	�]A��c��v�p>�&�7��Y�n�m��2��+��	�_�[��;;� �{���~�#˵�$�:�Kd)�:˚�o�<�։��e����aY��F��+��Őh>�M��'CCI�k���gvæ{4z4`y�;>�2�w����1�k�����h񜥐�.�n��ދ�ᇰ��NU_�$-r�����W�`����� �?�{I1G������Q;<���]����<��)�;�%%�;�2�w+�r�S�݁Cr����&>T�-dW�?�J.��S<Z�-�TN��@SE*�0�i�
��#w�,�7�k�l|-��ك����'s��K�Z���Eg�Ԃ�k����ݍ	�\q�/��✸�=ݮ/O��#fЦ�3?�\�Q�#��;_x����N!#����p%�J8�|S��.Ϧ��6�a�[;�}�YQuc��tb
���6g��M���x|�P�{�Vg�g��OqV�S�^I��bS��ž{m<�+|���l�ڕ�[ӬNF�_f�~�xg?����	M�0�V+P������s�82�l�#ʣ���pc}7iN�,�H]	sj?9�?��#y��Z;u>���ڞ��g+��^�ٓ���d�����ി���FP�2FE��')�.��ob�dqz�w���&�! �Q�}O̨�mz4y�7�Bo�;&Hǫ~������8��LF��&��/�X_��fy��q���̇�z���e_m���wd�0b��R��:E}�tt$ݲO�X}���,�'-X��1�L��t<ħ�jp\+PBm�l@i���mx��i��N���g�X�X�q��ΐ�<�1��;[w�X&�^M��ޕ�|��X���-1x�Է��oH��/�x���f��I�y%��/����!�d�@"���˝9l��9�b��V���Bc�m��e_t5�����@31:��Je�"WE`�b~;��:����ŶFh3{x����" ��rOG��Ԓ�=Eɐ�i_�߇V�k�����V�z��/"����5V�]�u�;��k^mw�+125�t���t��b��C�v;ПtE���d��G!1~�l"`x����`�ΛWz!7�O�v�0uH��yI�6��/�:t��"�k�{�SD(+:Ci�Q��iOZ�
}QwU��jM&�M���3׍.��B�3�^�X����^4�q�	Y	�LQ70��p���2��@��?D.�}pX�~��械��+(h�R[.^�C=�X��H��e߾�T矇&����&����;(g ����ј�3u��s�6�b�_R�t�	MY����f���$Λ}��(Zߌױ잶�o���3.�E|�X�c����Դ�>1��ZO��o��-Ӿ�:��x�?V�' �sb�7z��;�� �}ti?MRVىZ���y�}���:u|M�PO�fa� ]"+�Ԭ�ˮ��CwS�F�����g�ɽ����u��ݏƏ��]<�}�Y+Q�������C���q������C���}t�tj��S
~�uL�{�3Y	�O�}im����5������epّ������\����x:W����݆J���cw�S	�z۾���R�X^��}	K&v}��J?��y&��w����rтy���O��W��ߏ���&W��y�YB��I�l�V�>{]���z�g����t_�P�;ͫ���mU���6o6��⚭���0��+~/�	-=����CO��Rye�ݑ�/oP�E>�$''��9���yB�ϺRŔ������ĥCM|���u�M��vkL��Ϛ^'��*��4A[m������=��8��ўϴ��mh�կV����sJ��p��]_�9k�L����E�;��o�3�Q�
��eO$9b\
�m~B�]&�e]���\�[�/W!�a�%w=�˚�|p����P,����`���ozՕ^iQs��7�����L���*�T���7�B5:!V3��VCK��k���>t?�{>��erRT����&�$��͔g�v5����fa
q��v�����?����#�B��7��~�͡��#��k�\�t�g�B�����,�B�}䝹�_�h.�˿?�Ļxy�AP��[@���pz�Cc&0k7g�͟����ĭ�%i���;SʡCeR���L�J<��@5�Q�Ƶ���v��NM���g���L8��F��,qd��C=M��c��>>_)3��{������Z�YN��I��l�����d���ۚ-Nf��qj�ư/.��B��M�i��qnT���3��F��N�)��biÏ��E�KۻK;"��#q�_ym/�⯥��Y�VH���z:��u�Jy6F%�K�����%v�#'=,�3�Z��A�ܴXD[X6��L�D.�黨C����Ε�\����D.<��\4��!���xYt���|o��h���l5��9�%S�d�^�z�|6We@[��T�T�C-'�D�
Y& q�k}v���<z����[S���M��4���a0Qx{�ߵ�Kㄌ��C�,1���y��������y���q'�~����l7���y�T&(Ɠ�:��wyS�R�������SZ��.��	,�c~�����Ϧ�/Y:M�<&��M!(�S繻3�!Mv 5\��q{�o���&���Gj�f�
�1���Cbڃ�E��i~�^�_1�O��5?ʕ�eyB%����O�����U���+$m�ͥʹ�R��iv�Y�y��Z�$䚈Y���7!���r%���M�c}>I �������q����SB���+���N��s���d�e%�q�*���h�5?��v}b�޹�
�W%�<4z���o�aP�| z��S!K���_;ݜ����¦�v�~�� "�N�~2�UJl�6���I��\�u-�o�B=��dJ"��*2a�N^�lMSb����i�\��=��P��v_(d
?ԍ��q_����߁��U�I�<hB��GQ���Zj,�7NA��7�c��g�VN!�9]8�,���	(|B96����EA�n��X2���Q,H�[���@��Yz�$���l�Q�I�u���X�|�ԕx%Qq2\�eʽ�\p�)�V�6v�j�=����� r�th�td���M~�;�V���%j�L��c���&۝�a�`��=��A@�J㘮�v�BY�L-(~c\uFR�_��T9�z=������nt�5Hh���? @#kkc8���$Z��=�C�#�����T9Vz�Ɯz>@�[���U�����S���ܴ�S���Y&`��_g޺+�{�`S��(L�'�벊�:^Ylށ?#ZZp��	�03�\��.b��v},M�I.0E���Aw���լZ����L@��3���%.�m%#��(0+�O��]_y��f�n��֝�DU��On0N[��+�u��<��'��G+7�}N�l�:t�� ���< ��/����ئ�:q�E����G��48L��ؖ�L%���S�-�~)ޘ�������h���g��X�V��v�S�+�*���:���v�WWǣ[�yjVO��p4��0?�az(B��׭�B&Tm�� &Ţ!x��w	f�_�=����w�xC�F��*���{��SJe�B�g�-�n��z��(Wd��:���4.�jH���7��`�xF��t���
����������8qM*Q�@��7���׆T�B�W��������Ǜ�aĬS4�A����4�vu�}��9l���)&q��&����\���M��
� 2��1�I�{��@a�?x�'n 6�63j��f��@��)�f/��5h���<�X��:�{�b��L��Qv F��͒q�ӬZ��i�D5YJ;���>�̀b����^xS�e;��aeZ����߭4�g_����8W�Q'M���o'�/q��NOw���䒟�������r��w�����ǧ�"{�ӗ!C�Ɠ� ���'���ů�S	��i��/B�{05���/_T��1�U���;L�ofS��h�{�=sBd�F������]�㺂y�IO�F7nK�VnN���F*����ёu�n�<͏d���P
c���8�D�^E�X�A@u&��R�u=-P\��ڃҹ�����!hwpw��-�y����r���bo�"�wˍ�}(.O����.gT�����p"�&𻐝��O9����L~B)�@�aN�`,΄/nMFO0�LZ �ʫ��:�'�-��)G���;O���"+�[O����k��G{?�/p�E[�f�L��YǞ3,Ϛ%�{�|�b���N��5/��{�	���SAs�������ZK���`f&��U�W�J)����*�@Yg��$;&=̶5�q���ө.��[���8��w��t(��d��e�vd�Z݊�˨�bƖ� F�EE	 4(��3А��(��3�U��^R����b��E�V2Z�F�BS��`��	 �Eի�C�Q�d��C��w7��X"��!cX_��������Z:P�~qc� v3;��x�@ɑ_P�L&�wxZ����S԰v���D�5�-�>�ah�~���]*��Ʈ��&U�)���!VY^x���oYE[k;z�5z6�e�=�#ret��M��>�D�m�����iz�m}�����m��y�#���Gr \'E��y���l||`�������އ�8Ρ �����?}�#/I�ՏEkM�L��^�NU�f�yq�^w��V�`� ����+`I�l�<��]4j9��ّ� �&(_{i�"�/�{��ɷ'���I9�Q�/�������3㭶�l¿r-�Ô@4g^�}�x��>����6j�x�~�}ϼ�����>�a��� ��a@�S��g�%^d���'?����1>{��}+>����N�� -�EH.��{m�~X���sh����G�	`�Sβ���*��-������DFaJ(�˓��{��a����� �a�2�S�w�f�K7�(�5;٢W�=�z%�"c& or�w�?z�̑�f�����x�12��6����v�������X�[n��x����?��Tc�QGl�r�< }�	�)Z�{�j�-�%B�E���O�׿���R+8�OU�/��X�������ެ+@�ɚ�v�׉̶�Z�qd��<0��>Q����q���Q������)�
~|�MB}#?@� 2�,3iu�i����D x ��E_�sа���}{���V�����6�W��M�(�+��t٢d/��~Q�饠f�n�c�P58/�ҟ ���b]�T`��&�5Λ��E�0�-F?~BL����0�^�T��^�;T��	��������k�zW��&x2,�%
�,b��=��0k��
�a[��5^���nKfgU��.v�7���O�{�8vo��&���l�-�/�dϑQ�HEQ�>����N����G
}\%'�v0�PҾv8O_��$����'����8��ͣzQ<�8�rk"El�K�K+�35h����]l8Q�q��3��Pxw;,Ճ�Փ��0�iU��	GA�oMKu������#��-t�TO3ɴF�qɿ�p�#�a�{r�ki�P��니19�ա���)f��u�N7($C�ot��Ӻ}!��/]n���]���7N���Px�O���6/�n�۬��6%I撷A�[TT�(!Ç���5���Z��8�z,�My�涏�kڱW�8�7���f�#L��H)(�����)��.�5��W������z@�^�2�����HپokS-����Mޔ�L����8>�پ�┢�|�u���p�F�V���3z& ?�l�p��W��4 u�"�g=]�UC��ʑ#��+'V��P�9%�nG3���M���H[9v�-IQA�u��z.�@���M�v"�>ϟP�t{m��t���<�JjY���C�o��=�_���^:>��Z*_�ǯY���(�
�@��O ���e��#�+�m�C `d{3��n��$#�??ߺ�^&�F[�l'ۯ*�5����緸���sW{U��ms�c2������I�$��z��0�^X��7p&.�<Qrq�m��yJtu�d>��=M�joX	��2d�*������4����.���F�=E�8�����ol�}�u��2��hKf+�*�v�d���Á%����5�1��V{�������G�T��Ԃe���~���.�����m@�$t�����3�:�7.�a{��4��[�ѧ��<�&K_������a�2��ma��w����d0�ڎd�;�5`�{�h�xJ����������ahS�:�MUv8��.Yɠ�����Vv�0�kE[,l��Iֻ��naR�Z[+��k�*vk����">�ɾ�|����K%�&+V�C����0t��7��/30�O��(�~���eÐ�F�D�dћ9Li��Q���k�fX���|�C��"~��l��J$X���m���m��+7��i%�|i�mZ;��=Y�eA��0I�,4�W��<�AT�g��e�t��f;�o�`fj*�Ώ������SX|������b9���DT�!����E�`)&�0�>qw4���ڹ��YO��V{�,�s������zzz�8"�����x���"��3���1f�+�p���c�b�M���H���e�w2�RK��zK5">oFmF6��6W�ϔd�|"N"��������m��IgR�zim$�4>˧M%�+�]0��ׯ�4KL3�y�M$f�4�����H���CKO0Jw�D��9��|'a"�����ǧ[�nwO~(��?�|��b ƷF�D�.��ӫz���	"��&8�)ߊ�e��"�\���L��VyI{xz��nX�>���B�.��9P,TCZ�g������n�Xש///��K��� ��G@�&)�MKdR��FI����I5{1'������N5�V��~c镜ʪm�5ȧt��X>��s��R��;ZC�	=^��F@Ʌ������Έ,j�����N{�˓/Y�v���ݛ�7����+'���x�����&�IN�I$��+�Q~�X�5d�絀|���g'�*u�@��k�C^��:����9;����RT�]T�8��S�@�P5���JY���EW9(��ltEl������w�"���6Z[+����=�Ӽ;�����\ZZ�5�);��_Z1$�q�BP@J��-=2��k~|���m~�b������ԥ6�V	���/�Q�9z�w��y���ȏ��� U�W_O��T�r��x��>2��[r)'k�z좧\��Л��?��J� o�jн��a𞦆"����@\��m[u'V���L��?�gv|�OSy#�b�<�Un":n�RNx����Zn��M��n��+�����I����Le�5d�H�e��)�#_����tA�j��C�S�g�O�7N� �^�8���x�6i'á9ᙼҫh��]���MvN����񙟵�ݍ�'���,eQ���!��3��0֛��vO�Z�@GMk�m���ͼ��4]p��Uװ�z�r�l��b���H���W��tp��<V��Y3�Gz��>��"�g���n��չ�O�Y|�!���u�q-�I#����)O� ���c�m��� �஍���{�a��M�%��UGw4�(5�;F[�>,ׇ�
f������x��3˽�w�|��,��쁁�-/ӻ�Lxə�P�nk��Q��)&�x���}lt���u�Z��wh&�5?=�<w�2r��9���%g�� D$~w��ہ�Ĵ����ˤA�cΣ&V���A��p��0��Wg]���)��C.3V�.[-.��I�^hPwG�a�
��!I����OETD/[���۝T�*_i���.S)Vl�{1�x9r}���U	��XEc<_#�@"1��K��� i�h������=��n�r.|g�����͏�fVOZ,	_���a�8	#������	N�S�h���4�4�5�X~���Wf�us{���X]9�8�/�̐!q�S�|/I�����Z�T�����h�7KK�:�����'�^kC�ܭ7�$�W<ȭ� '-���(��0������VC�!���pxt���Z���QÀ�a5(���V��G�������!��'=N(V��Ƕ��ZK����w3�@�G�����; ��TX�w�<>��z���dk\��Z3�54��vm����Vzޖ��JX�Nq	������<�S�%z�$i��!��̱���_�&��]C ����`��I�0C�/}W�B���o��2*eD��.Ɏ%��N��i���]�� _�N�\��eU(���J�jA�u0�����\ɮIB%�*^To��8u�$�1�0���_�>��}�vQ���h���k��� 
_�2Lx��}YR���`%3���c�&�oO���sٰ8�j��ñ,}�}X\�J��F����(H͚Q�������ћ7N�|Z��(�s�U�����gC�HC�����.����!��$m����Z3|Q���f�}빏�	Cq���;֢���ᙩߒr9�f�P�
� �����?�hL�-�MP�����n%��?�!�6�z!oKI�c�����W����W&�����V::R�d#��&��2ք&�y�N�a��M�f��`г����T-t�ɠ�JE��jOx�j����@��U��8'��y{^��0E�PP�%>OJ9Oar@�{C&lB*앧s�s�;��R@;h8l��M��0����{��T綕N�g�(M��}�?��p&,��	��6������'��xs&�/{��}��D
9�	����� QU&b������e�<#�II�|�_&���&�b����L�V�X ��W��L���M@�F����f.�G��:�}�Zv��M(*$
z�R3rƤA����jWD.�v�gh���Ӱ͡*�~I����̪�y獵��0%���W1%Z�a�Oh��?í����S��O[o��f�?&&���+FE���RwMW�� H��݃���ھ˭�X$$������@S�Q�T�[��d=�
r���~A��v�p�ɌP��ȕ� J�L���O���)��"�쏺8�V����fI���G�Mp;�ؒ�d�ꔷZ�rĻ%����ϐ
�'G%ך-WqE��#z��j��ˉ �Q���~��cF���f����i��^x?�߻���o��?a�������rw�^�3�i�[[}��[���UKF���l���NcZ���	%�la21�"��N�o��?�[����@�1!u���?^��q_�/ì��]u�mB��æ�T>�B���G)�j��Z3�F�(x¥��?�p�c;�߯5��s��_�VY�[@�+Ia�rJH  H歸�S*"� 幢:��޺�e�V6���ڐ������[��|؈D?�@�{¹.N
1I�Tqvm�'�1�������N����C%a��R�:��K9I95�+�NYf�*�P6C�`�BEYY���RGXY	.�)��k� ���{��l�t{"�������I���Z��Y5��P/�G���������es|����^;kȪ�{�ldV�74�:�r�ev�
9�h,շ������4^_����_=n	̕�go�"j�5��,"��K@��y��)/ΦKPy����T["�����9n��R����YF,,�մ(:�p
2��@���B�nƟ9�n�ҟ���co9���[/���&416�t�c"�|o������5�0��.�V.�)*2s���3J�"%��ڨu����v�V������JJJ���l�����Bi1�-֫5Nj��j��L0��僾�9u�i%.�1.iڃ�+ŏ���3���u���>���3+?���tS	|�2��À���g(�=ӌQ����V�6�J_�-m`���l;�~�z��W�d��g�cy��V���B5��S�J�&��o����A����b(�Xc��c�3��􂞮&��-��3Y2V�51�B�����h��2���Do)����̎R%&{�)��!ފ_Q/����F�|ؖ��iLy�g��W^9�1�d��� Ј0�A!�wbT��^��x.��}9�54q|�� �a�g�_9�Lg��-��hp���e�ti����`�IUZ�@��!�u�;�E�6!+���͋dxє�G���r�"T���Ă����P�fht|�b��l�Ą�z"�����Q�>9u�$������N�6;����ٿ��ȋL�F�D���)B�J����̋�o�O5�R����݆��4}��ob4�Jt�Q��S8!=$�=:�&/"�P����T���>̵�3|_�?�OP�S�4�P�,+ ��=�	ϟ�H<3nD�EϰӍ�}#�#��cs6�AѤ�1�a��>���V�&�p��:q}'C��jE���֞gw��.��J���%%�-.θ��ڞ柲�2e~�m5�5�3���'�t=��Gٮ����U.}Ň�̟�P������#t��N��L5PGů��*���]�H�ؘ0V����5���ͱ�Y��M	�RAF�7,l���Bv�H4���S'��VA�<ڞ�"L�S�'��k���M���ۈ�:�0����q��ث��;9�"(�x^b��;Ze���[�&�`��-�5F�:�U��* ;������O{ʱ��6����6=9k�\ﻹ>��䍡�Gb����fT�s�)�V���_�E�r���@|�=G��J�p�O�,?*ڪZ��x���?��	��LQѹS��v��V7�#ug@9���_W߷�~��6��<�&)��y�;����|c��� ���a������$^N�F�^��Rkk�D���9�N6����M�x���E
��ᄹV|}sssM���Q���9��U���Ц�Ͽ1?E͈��]�ʉ���ڷ�e�V ��Ӛ �Bd��R��-O���� �ɥ�\��6��QI�����M�u��j�PX�^��Ò>%�K���Vm�k�S�4ެ
�?��]k>Lָ[�L` HY��ɼ�����j�ޮ.?�H�Y��v��g�]BI��#˗��~]��l���>���5�p��/��@ -L�4�m��m�.�K$�m~��\���[5J+�.��F�X*��jd�J ww�ܚ�ZO��M�ȏ��oy?�;����׬�.L�,1hX��{��3Y�T�ɰ�1�^i˰�1��7��[�㮤����$���~��*I��6R��D�B�#�H,�SJG$���S��D��E��h�Wș�@t��@n?�h�")��<C^H�6щm�W�C��u��8�2��x����^wP�]h�:�������C��w��
x	6!�UTi�	�1ԷW{q*a9�J��=O�GhCQ��N��yk�����^�RRR��S&�ͮv�m�g���ْ2�)����E�#�$�G���j ���d�5����. �W�1�O�*�z|��h��r<�"�L�[�x��Դi6=+�	1]&G��K�N�`#3!��q�{IZo��1�����,aBҋ+^]VI���P����{�H�q� �r�8�$ܧ~�6,	Y�Z(-�a�p��HsN�/��������h+6r���%�*�`
�u��×�II���e�����K�?���nr?S��ٮ��	i�ME5�A̓�&^f3&|n�o9�U�T�=p� �a��!��Y�&�� �Đ�6d͝><��z�x��p^��+O��l�oF�:A=ż�<��txG�T�[��3@���U����yV'��aBQG��`����8&�:������a:&�JL��&{�[��a�0N:��총��Ĭ8sZ�%cԶ�C�\P��K���|N�T��Q����l(VƱa�q�P�6�z��r��;�m$�d��r�ÒU79Q1�ݙ��?�o����q-.2딒��%��z�����0�-gef3��%��If��&R��Rɜ{�斮�$�(ޢ�pKM+%4ˉ��ix�Оļ� �Cm�缻'��G�����������8�9?C�٨���H��������@[���t��9lK�������>��\������p��7E%�hKoF����L�����bS�-��G���-ؙ4[0*��]!l�%�O�6�r�Ϛ0�W����"��H|"l�jN|3U�����Uw&�+gf �*�:�7ӼiK�@���A�F��/�oW
M4!sCa�m�H�l_}TTj(n�C�^�)v�޺\�����eJ9ͥb0�u<����7ip�]�Pr��!��v�%�g��]�E���m�ct�����Y���������9eEv�,ڛKE$�ħľ���aW�gC���X�׮�<mG;*���E���'���9x�N˦�GMx��������,T��Q���"���m�%���up�言Iv��y\���΂�68�Z�k��׿|�o�� ����~I.�W|U��*5����C֦ӕ)�;�V���Yϱ�Z2h���Y'!�i���Q�a`�?Juf�+�M��1{�O�u����c�N%�z��S��B�x�Š����b�q�j%�����0\��[!DG�Q]J���(Nd��l���'�{9���p�J3����.����ϙP�ut��ߧ�����Jv��^�qw}�re�~(����I=o� ?5��J:?Pj�GP�g�5�����z�H-�q�a�b���<d���2ik�ɋ�c�sZ��M`Ë��j?=���PIb��r�Gݛa��Wj��-x�p&��G�K��7 �p7�;�Vg���3�i�9��R� J�������U0c]$U[e*�_Ɲ��E���CY�q�$�nu�l����Ŭ���p���ME8� �g�	M��^������1V�+�l<1nb���%j���Ғ��dѰ9ٖI0�c�A��ToƷo��v"�J&���,��<��4|=߳�d` �l���@"Ʈ}�:���o�Ò���"�s0F�w	�??έ��!��*�1��t-8�p�Ԯ�S;�e:9>wV]�L����F<���ӳO�����*"�歙��_��_�V����`� �ݞ?�3(��X̂�!��y<ܒ�$�v��J���E���<��i�M��{z�a�T��(yr�v
���C�0��M�/��x�;��PK   �p�X�J �i P /   images/6a99ea4b-7804-4d0b-a50c-ccb121b20ed8.png *@տ�PNG

   IHDR   �  �   �$   sRGB ���   gAMA  ���a   	pHYs  �  ��o�d  ��IDATx^���e�q�	�u��z�M�n��4� 
;Z��ӎ��w$�ҎF�!5����5II�FԌF+CI�4R� 	C�h����.�e���{���8q�y�^ջ�]� ADU�sn���Ȉ���<y�I߅��w��]�.|�߅�x(d�o[�v�#gϞ)��%� P2;Z&����/��y��k�q9;�����y���ى`O�� �ᜎ�BZ_�G�Z�g �7Н�Nօb+��;��t`&#=Î�����(`P�p�����j�++�]�b�ĽG�ΖRiR�G��r��)w��Nэ��.t��b���#A��n�r�E;��N��h2;�\�,��&�(ǎ��c�����o��R�C����N���RA�BQ<v��[GEeQ�!�@*�\���/�b�5�:�<;��նv��muş��Rb�THM5��ju���Z���#�����oZ�\��o;��2�������F��F���N�yk!tSgZ��*KE(J�J(
('���2h���l�~�?H1[~� �4�7i����F�������?����(����28]/�O�,`t=��z���Y����RjwZr��o��R�\8Q,��Q.��y���ψv�I~����V��6vf�̡������'��P��]����-��򚒰;~o��h;�V:�=������o�ns[�.�]����4;m�}�t�ِ'^n����T�_���݅��'fg�,Z�o��[����M�Z�O�;�OH�7hH���V���!�R4��1r].�oCB^������5�n�}�z��y�m�:4����Gݔ�E��:�3F�mu�W5F|�T.���������v�� .���۵n�ժ��n}���w�RH����wO��1�>h|=���]m��'~_����������߫'��)��k�����e�����|�4:�ϧ��~�޽��C�t�''ΝK�6����j5>��堧�w�p����߃J ����^��
��zԑ�k�:H��7�H�7�<��t�e�i�5m�#@�h�žʣ	
����GFGijj��8빾u�ӈuU@�,-o�7��n}L�2���`�<����b|g����KѹԵ<��;��y"l��nw��l�ssc��U����p�.~�[b|���ex�0�	�4ó: \�y�\���3��iyd8��vy�Oy�瑾�����0�?��FZ 0�6���L<�J4$5��fЙ�tZ�V�^_�QeY=��A_�o���.T���7k����v	m,/t�Ȓ���S<P�S���f`¾�`�� ol�c�Y&�'Ǹm�.v-O;?��q�r��A�1�3ZŒ�gS�>A�NP,U^,�K�����x�ȑ��[ �� �UΝ;wg�Y��Z�^ocC�+�����}o6�0h$�|��B���Ac����(�;����y���,VG&���|��Nc"֧���#.����luS��iubb�禦��=x��fV����媀f�{������wI�s���Oao�Ȇ1j�v�+̧Ű�-��e!��6�)[����������uأq�6:nM7Ϧ�m�ua�����B�8��V�q{���=�Ri�U�-�7��$��n�yS����~�����F�6[� �LJ1D<�y;��(M�R�y�\J�P]��H�m�nKu�,�����R*�E��T�RɎ �A�R}]�!C]ku�J���X���V���;gʈg.�Hŧ��+�_I��Ie;�g�v�B��B?�pvOg7��w����g2"rA����T;�v^�5�s;��J�;��G�K��9sf���}O}�A����յ�J��G$�C6ܪg���a	�{C��4!�|�'�b��X��>l��P.O���Pl�R�߭���R�O�|��j�i�Z�6;g��s�RqI�6�FƸW<�)d��w��wJ�)�ʨ�!�,D0C�7�]�d ��|�whH�-�˝	$Ҩ/���J�#���n��������-�����J�Ǝ�?��{���OJ��፶�M�)"P��ƷU�}�*|L��*�2g��t���_Hj�e����f�ͬ7��Y�ח��T,��)czd�\yn�R:7R��(���Z��rY��z���ڬ��j����v��2�I:Y9361T�`d���x�:$i����v�O��c��A#F��W*=<1;�w���~naaa5�����\]XZZ��ը��V��#���͆�é �9�p���u^h|���tYC�	5+�7lһ"�E���y'�G|vXo5��??R�|�T���x�陙�ř��F�p�7�UVD���9ӜY_o^S]__�Q���n]�])��ʒ�
1���9�'�/��o�$����9���%����yytb��/���{��L����&��<yr�R)���h��N��>	ܼ�����BA珄8y!����u���b��D�t$��]�(��a����_����]?s9�A�/�}��=K���77�?��OƷO���np�ǧ���q�o����Q �`�����������,�*c���M��������[�2_u�7W	&&J�����v۷�p�Ƃ&|I1o�p0����c�dF7�~a�Njh���ȣavU�o��O�o��ׁ^��e)�����{����Iџ���D=ah � �����y�������As��9�N��F��}��s�,���j|���|�f��W���oL2��ыuёs	%����B�SR�Fa\�c�7Qy���}!*?ld���j��ybjr�_��-|n��׷�c~����cӏ�OL��8X�7�'��e��Ч���Ʊ��-�v�Q���a�0\v��;W�P#�~K��u�&'����3[�o�c�Z�my��y����U5�����f���-Rl%�|^���P�`���vy�Z�<�۱�Jf�B��q�.���kf�KW�����/OLL?R.>�Iș0�>?}���,\����,:���v��ٟm���#�j�}����,��U3��������;��G?����Rq b��+ �g��=a^��]�f�Y9��!ʄ�Co`�Q]j���N�N����ïf��>|��b��h��x���)�p�>�����ImD�	�PF�ǎ�X��f����w��g����V���μk;�j�v�7��woV�tߠu�����HpL��Y�*E��cC(�סּۥ��,7X7�Z�&ٷ_��������K��gWD�9==v�R�|��n/R/��{�<OW��K��c�,��~]�^}�J��.�W��������Ɲ��y�k�oih������6)4_�	(0�>*�iZ:y)�0��;�K�f���U*�o��=w���y���p�P��&����C�)\^	����c�hy�q��ah��>F�AD ��P��B�V��������Kcv�*�U1�J�{���|���^�g������b@>-�����>��@�{䍪�r����[b(���F�N��Ӫ�?ֆ����6�c��>o���SȂ��)�� 7�W�޿xr�{�+n|l�j�[�(6y���=j��p��5�B1J&e�H���d?{�=K��#4�F��t�����+�s���
H����,+�Ո����6�7�|p�"OX�����f���94l�U.}��4���2b�Ni����Bc���Zm�M��q+v����Z�v74�OJ���@��r�H��<Ƶ�֎�/��Ǽ��w��B��_.�6b�*�J0U���˥u]������|�L�a�5/�' �y��������FY���k�+^>]ޗ�*pE�osss_��|W�Y���jL�07 G0�Y���ѓ]8x\( G�ؚ��Vc�o0=�����o4��N�PCW:c�b��*�b|�o^�ls��ہ��(`xH�6����呌����|�ˆS�}ǚ(�BN�Č� ��Uݬ~hcs�ƫ�]1�RG�����V��V�y;S�{�h(�b�7� ϽA�?���B��|����s,�Td	�R�[�W�me�
�v$(���l���8�/���]��!�A �zB���y�P��k�T��x��b媭�]1�///�����ݡ6�橁�t�e|�8�]��	A��-�����	0�����e3[!���&ʈ�[�FxR�(Ք��R�eyn���0Z(w���G�������T��.���.�L�aP��E|�'���s�{F��M�(��2�`/Dl�#�9s��sζ1������F+aj�����/+�;vub�+b|¸��Mb�����t��{)���e����\�q�n�[��ZGD�c(��^�G>�+�JJ��½k��j^��@�ژU�Z�i���V4:x��m ���o�\ۤg�/v�4��]X##q3��-��h��Qk��T�k�0\�[YY�߬7��m�ޤ�4���	T��@~Q��0��(�9z����øó�X�������B�ߙF�%uy��f����f�֯�<At+�k+��u�B��ݞ����Ӂ��0Ѿ����Qli:�l�݊EvO�5IJNC9�:�S��6���z��=k�|O����u[`bqS��������З�у��y��"���7*h�!���,-C3�1d���|=�3�nwn�7������9�+�ν���^�>�R{���cZ��m`K���q�JA�U4�ͧe#r�d�sy��-Ս��.���{��W_]=� �����C�+�'fb�j�K�p��4�g�!��2�Y�S���JӱG��	u�㉰�gw�{�x�a2^P<o)�n�@U~Om��޵��(��ID��x��M�z��bi�vg��JI�'{�)��Y(�o��j��r�@_2��7$j�#�|��n?��:=��2�HF���/��U��د��fm�MW�Y��%�n��T��x����X�G��y������<xZ�@�4�n��(J�-�.���Q�փ�s=��|��\������Nx���+������]Y^��f�6�	#-Fud���b����Ӡ��0�0��Ҝ��߲;����ʍF�͍��\�'�^���[��ʋ���{o �kMy��Qލ�zz@���E۽%����+h��t�x����V�ul�j׬�����ųZ[;uEn-;�̡��^��V���r����ldC���ډ!�1J�>�e�	-�@^_��.���l�@FŘ�B��!�!'Յ�8�:�&��oT?���y������l|��:�M�!�����v���)q�_�����~���m�$� ����
�}^HC�\G��V/k����,���gO/~h}}�u��;v�����]���aq}m�R.�h#u!x��
�q1ȷg{���˧��r���ѕ{E���ʹ�T^�����l�o��o~�ө �J�k6>)�<�����%<�z���|$L�Jc�0B@�\�(��?��`��t䶇�s�z�.�=���ut��e�RaD�UI��g/75>*%� Q�z�H��F+�V�u���s�������Go���>gn .z��go=w�ğZ[Y�����m�g�Ր��&<��\`�!"�C.`�� �?3Ҹ��=ϫ6��f�$Q��Y_%��0��[�̮Z��յwhbvE�����L:��U,��z�mD�Ʒ���'����	�!��=>n�D�]�0�	ф00<ش�UR�z�B(�?����YqM�,@�/4�.������5�B�o{J�������s�_������S��SS��T�!�^�@��Ley�前��޵͵[�7��okkk�[��K�گ�׆w<-!	i[:ں���_��?��v���10��䤿!�8@�{�/��3X��Y=�\3��Uetlujj�w�w�����+��ڌ�5_&��-޾����n��'���b:d�ftH����z�r��X�`F�-� 	���AB��a�J �i�}�S���ə������dQ�V6~Z���}�r�bˣ̥����������FǾ11>��he���{��)6��F���V���l�V�v����F�~W�ݺ^C�.4oW������k#e�'ۅ�v3��S���m�c�C;x�B\�ne��r09g�ށ��$�]���|�#���{Q���g$��M<7?��s���y�u�d�B�w 1>%��)�o�V�m2�"�����g�ʌO?�FΪ�yB�0>��!� +�?���a|:?��2���ax^�+�s3@y6;�.�,?�e�7o.@�q�^��G�ľ�b��2:2�Z*�7��b��jj�,��
i������f��¤h�b��z��������Ė��:1�P<�ubǞf��:����h!O ��h8�|LȀ���o�lD��U*�:J�������Ѩ��������]��P�-߸���o�Ɵk7�{-h���iΆ[Ʌ��oٹ�,��	��근���ڤB׹�ke`���:�Q��N�3:T0�g�'ۭ���/���<%��f&/���@�GЪ�<@�(ó���%��:�kf��lW�"u����O`|�#Dq޽^ o|�?��AA�Xݙ�CZތ_�� h�o�F�娺��8w&7zh�<J h򜚞}ezz��.,�sss/X�� }n� 1;��|�=�Z��;��4kՒݧdX����P��
�<ݮ�w&SDN#f����P��r���ȉFI)��bb���j�53F����C^I�)So�8�CHiQ6�s�p~l)G��0B�#Bh5u��W��Ŏ�̮ѣ9����|�Fm�	�d�����eс�7�4~���(/������� �fm����ع���:����B�+��!u�������c{�������ggff^��r|	��8{`uU���Q1{�����1��7����y�h�ݓ4Ad����<�� p�C�а!���f�\_Nk�,�b�c�%��������&ifz.�OM��I�6��[��ѧ&�-ؚ��!
��*kvnl-�'itr*M�L+8��������༩�d}e5U7�Ec�h�*?���Z�,e�<irr�Bx�v��r�ae���8nɃ���kvn��a��c��ח��F�Ά}���o�ͫ�v}ff~����3��Ѥ˂>7C��ҙ�7�k��n}B��4[�i�5LB����[� �^��t���ɸ�[��@��ѫ}��D�ܮ�\�;R���sieiI�����R�3���-�KD�g/(UCE��`ZXX0Z�j1�n���tӱ�G���J�X]S� �V��T�њsRm*צ]2�م�iρ�ifnV��p]��]�P��L��ϦWO�P�Y3ZS2,���ƻ�%9)�26����g�l�=e`�D�����auY�:��gymv�J����2�`'�v���f��F���y�r�^x{��s��4�����ߖ9��F�,�`TǸni�AZ��c�*�T��V.8D	9: �nuc-�;}&�d���b
T�F�a��I߻o��iy������q���RZY^J���ehM[���7ާӔ��>���B�����;����m��-X�d4�[�71d<�����Eձ�
,�([���GY{��7�v�8�c��Q�v�yI6�j>'Yy�	#�a���Ǽ� �%?���N����L��eet�jw[j�3������s�aH�Q�4��MM�ݛ���n���P9��x)���5��f��#��Q���K����WFd`��s���|*JW <6*E�Ɩ�����Vd4�k�7օ����i�W<k�R�a�x����(1�.�ڈN f���Z-5��T߬���bm��C3Y�Ic�1k׈�7b�0^���F	�:��+!l�X����# K�����q�1��M����?��ˬ��3�Q���.�H�cv,if�L@[�S���Ïdø|Dq��M.�!ah�k�Z���Q%�4�ʌ,o�q�kQ�G�� �qY>Ԏ*k׳:��S��и��uks}5m�&k+2>����e|�:߬*6�0Ȍ��=��XQS.z�@���e\Ķ5�UOX�������F�}&[�FC�*24h�T�Ԍ�թs�_�Mʯ�s��?xT�a(^�XI��f��6�mx�Q:$E.������2"�:�����~��)��f�7�J2(M�z�N�,�8z�(�Q�mܭN~�����2��I	v�*1�
H J�I����Z�:e�.-�:º�(�6(�٬k�Ï�R�Y��ڴWS�����s��"c��ȸ�4�K�Dd�A�k6����U�uT]>T/)����Q���bTT�q$`m���:v�͌����9��:˦&%��ֆ��Q�<�u�N�����;��j�>�������T���t�d����J��y��T騼͔zm�f>6�P�lk����A�sa�df����\GK��fQ;1�դ��c���T6_�dx��WF����LPx��o����غ]�ƀd8�����<@(+�M���#�F^�_�)3ȶ��N�n�)�g��s�j���ڑSe��C�#/�p��x���E�X;g��7ƥ�ɦpn�y� 3�R'}�:�z��P�'�~qTL��+G�`� 3S�c���ye�hd���q�^���#��{�f$�p(�(��0U7^J�D�m*A�0�x$�Σm��r�W�����7�ɳ��U��b�y[�?ꉶs��"��6b���ݼ��)��s��0~��S\7YQo$m;��kypc۞��hK�Kj�E9���6��FC��\(��Tׄ*,T��<�	��[a	�2�TF�y/���2��Hv�N4��&�	Qv9��3�ҳ1>� ���dƆ��nfX����~@</ƠsLc��}c��� ���͹���E���f��N�w��m!_�2b�:4D�n�C~�F �+���Ґs�Ax9�G̜Id��� t	��%���C?盫�Pj�;{���H�zi�h�<�Z^_Iy��PfK�*I{#*4�����}Z�9eLA��$pL4�c��U3���u��\�k�e�Pą�A 墍����xf�s��]wT]v�E���P*h���4b�4�r͟��bЯ{+��DZ�j�o9�¬��GC�h�Th�g�P���H�-�'ы%6C�h�EJG�Ub�� @}[�i�aP���RZ>�h�3���E�C�R��s����%�o�5��RG�{5=�^��"^��-f����bG�s[��\�'��~���-&�H5Ѓg�<K�����נS�L痜w�ĵ3gΤ�bJ�Eu���6=yP���ty+���L^qD��Qv��v��>0��zQ����5�Q��ꊈ_�	`(0�t����;ߣByT��ht`,Ap�Z��W_}5=z4�8q����ϧS�N��"3F�P*0�|�<�X�.Z�x�Cѭ�q�ܹ���W�/��^y�t��1�=�N�:��?�������mkr��^Q�!�Y�Ǆ��h�WϝM�?�Bz�ӓO>�>��s���^NϽ�bz��ұ�'y<���L�Zg�?�c�� ��ρ�~��u�,TTW��`X���)H6����.3��p�S�J�Ӊ�p�����7ձ�����Ԍ��V�ZO�k������aX���f3mn�F�٣�-�166f� �ESã�`��s�B/���F�W�ܬ���ʹ���6�{��h�1�MVx�M�Q���%(��V�H�u&/LdTuG\��i}C�ա�75�CD��@���k}�D=�A�x������c.�va�E`X�c��f1/�p�0��y`]� �!X��-�f�X ���pH=��؄�q2U�Ħ�"^:�K�77�0��53EWk�E��Qgy����X�
-4V�p��dȵ6ґ��v7C��3y4^�����X�5�+#i|j*���b8ޓ�ԐYV[*��i|b&MMϤ���!��!��bx� dC=юa ��"=�c44��B�ex�¤�Wh+��[��8R��q�x^`2�#��
�a)��q�FBB�e���7M�3��ܖbl4��L((��X�A�r�A3b .4����ǾP�o���f�y�����PA<�ٷ=_"4�W�a������Q_�&f����l���U�Q�W��#��z�i��-�JO�L�,4�ę���%������v�2����<�$+K��\m	�:��r��C�b�15|�N�/4���3�7��,p��
�{���A����w���C���o 8���ѣ�5\.�0Ɛj�+�c�ME�(����2�C�[Yqst�4y:�s����!��ȍVӼbm^F+
�~���L'N�1O8!#���5�����1hv�q�Ao;9�u ����� MG����f�`t���$f���ƞR�3ߐ`&�*/oh`��FG�2d���sҸ�Cb+�.
�׹O����}2��4>6�x��^x����O� ϩ�9��փ}��FZ��0�;�E�����M���]Q�b��Ȉxq;y1؏�O�UņO>�L���4�x!U�NMΥ��y3p6W`��O���/-AϮ�|2=������A�fV�V]��z>)�ohL�����4�3��Ȳ4��`^���!��D�`��Ɇv�Z�ǲ�?��hT��(e�iU��W��HO<���Ǖ��1a�,�")�	��s�d��C*�XJu��C�{�1�*ڵ���E��zx��?��;)j#�I��N�S��W�7y$=����F5�d�<ܬ�A��M�IB6�*�f�m0�bh���� �o��}�N���o�Q�tt#1�f�D�%�a���#�_{z�s�%�^`�6�vz�g���9V��jL �*'gf���]ilz*UۍN��^G���;��r��ַܙ�ւ|�֮h��̲A�e�k������������`fn����6��W}�J��!���`�m�s��U��"o��;cZ��Ď�1��{מ=��׊��Ç�I�H���B�	�E�H̘�ك��e6��{l�kFo�P��j�ntջ������O��_�4@sGX__���j���L��
l1,�����6�z�%�~���Zh9��G���NR���6d$�.�X߰�Ilxc3ժu�.���o���k�^���1sdd����Lyږ�Χ�gN�v'���
����w����܀߳����0��d(~�.�bk��s�geq��!YP��g޿�Ś�v�2�ȓ����oj;�	/��d!H�`P�
!Wxw�K�� �1r L����������*^�؅���%@�w��o	?���Ӆ�7����p�4*��%�����9#��Q^�0~�������J�(3�&�D�-�H>��E#>k�,����þ�-u��#�9�uy� ��1T�����4<�=��b,�0�n��'����g��Q ��B��� 9���30�jy�s �T���F�y�L�[`@�ޞ������s��2��U�fX-d�p���p!^
zy�y�lW��43	��^��o���*+e�����es�-QpΌ��,w���1��⋶o"�a��<����l����9-����3n��U�i��� ��=�aܜ�?�KCiC/�7��v�(>"dw5i� �v@�q��z��F��>C;���OM
��-�0�A��y�C��� �9��~�T˥���5�#/��BYS��¬sd��P��-Բ�Gh+�(�{�d++��e�2����Թ<���Q��=�Ƀ��F���t*�'�$dy_}T�.!��ѼN�9�j�-�ӹ4���Fڬ1�����+ă���N�G�nb>���G04���?y^�\���������	;���]���P�0�; �!�{Xo�ֺ�b�P���`<R$��rk���d�w!�]"~
����^ݢc��xTiʶq�(��0����8��1KF׎ޡ����e�z�H'��4��������3�v�MT �҇�ȟ�{= �<��^\��!<F^lЋ��@��1�u����D��9*-�,��˖.b�<���,�n�)�ØFku���?a�^:�ڳ��^�[kB�ed��H��"�.ވK>�_AC����O��,�#����uJ�Q�l�[6�aF�R�v�eBN�{�8� �.�5a������0��2��Az���~�� �l���p�6���@�s %��gO,�qh"M�o5�	^&��J�Ly����Ϣ�3'��`��y�Ǎ��X��3�+3f��mB�4 ��7�����lA��.h�!�Y�z�s��lW&�y�o���m�;��d������B(�By�� 7F�>p-SNV>� y���(�c!U� ����:��ZC�{,5S����2e?���2��*>�;���CRr�c<�x�(��QO��om񙕅N�:�@�|�]�ߞ�i�-6�T��]V����x���i�6ႜG�9�����͑:�	�,Ă�� �P`U� .�,o�1�P@�y�x1 ����y%�-u�fgm�\`f�4�Xr`<�P��C3�Dd�Ύ�	���)ʕò�v���6p�t /��q)Z@\�:F��|`���?N@/8c|����N�	!Ȝ���y�4��ը��(E�b]��Z���X��v��G�f��F8�E������-گ'��j��<�o���G:��]��O[䴳��H���n�:����^�V0�dG��z{����N�ٓ\����!���Zlk>�,^�1>Ջ���c�_�!q�2���8X.����i�hC(s��s��ᅿs����\�c��|y9_dΰ�RO������I�0���G��s�N[h|g��Г�hF�c��A�S��% �/��z�;��_`���vg�_l��Ł`Rule ��`z/���a�\���h���۹b���G�1h��f�Wh����X��Y�~��Ӷ�,U�1ڑ��"���P1fQs�K)�'C��Z����a��2D�����|	Æ�(��L��t�"?
����Ʈʃq���{"m�1;�XF�� ��9��[�;���2^������ v/	�
�]B�y����1#4P�&������8�|M��i�R��,���mk��<��8J
�	ڑ2�A�J��1�n�wų������Yn1�A��V��73l��BB��f/HŔ��?R�߂3œw8��������,�x>�������q};��-�O�ݣc��giԾ�����(�Wʻ�.N���2�k���>)bel�L��#�P��^A�0~��3����~�A��!��H��z}L�ӧM9)��-:f�7�<��qn�ˌ�3ڙ�Q���� �^��>U|���B�>��t��)�it�`�s���0zB@�6��������~���Z�i�@���y8��Q6ʓi y,_fx�?��~y||��OLL��ʭ؅�K_h����b�I0Ø�J`�kX*��� �w�#��P8�$E�(����]&~��H�F�z�d�0�M���f��˒��o�7H?���6�ijC���J�*�����+�'G��ky��H�R��A��a��u9Q�D�i�c��o&#;������W��!4�����İ�->^f�G��:z����,@.*g|��ܲɴ�3�9������n�B��z�*�PÈ=s+�(F+�Y3E���L�ƣ��d�c�+�b�҈��.V�u�t�u<�	�=O|����J*��~�ƀ�F����m(����kUD���9ڱT��Q�����1�^o+F�^Ӧ��T[
��=収���zb�;�mci����kw�`��xؼ,z�7��?o@��J%��=m�#��t�mk��e��F蚧�q��M���M�Uݒ9��]@d�N�`k�6�R�[��Ꞓ��S�N��Gn�n@67MG扅��/��������o�'>�# �KBf|w5��ow��˲$(	������4Rm}5�y�D�X[��ǳ]��0�Ch����4�]Hcxl?t�1fÏmQb��0��>݆�a����|.�>y,�o,����ߴ�Ù�߄��s��5Gn��FR���k�h�ІP��Ǳ2RJ�K�j�i[�9"�fE���(�z�����k����q��� <
I>���n*�ȇm���zZ�œ(^ސ�p����c|������쮆6iKe{������U�_S=m���e�7V.��2a�ᙡgzm�-�a�8󛇮X����[~�~fu^�F9`ss�O$�O���Es�aw���׫��h�ޭ�ev���&�S�h5������JQ'�7�6��a��)�.�Y���TUY�F�P�f����=������CG�7�Q���k��Ui⨑
QVK�����ڽ����GG�He�~����R$�����L�z�{��Ԃ�D�xS�����c��iXy�GD�����m����H�}��Y6�y����o�-WͶB�E����0���_��_O�<����`R4&1 ��NOO�����ZH�^Sڷ������5d�q�VdKy�r�̩t��+v��m&ބ� ��&�H333��N�>mݯ���Ca$�A��ɉt��a�;MN̦)�����>I��V���]�?599���k�*��/?�S?U�tը�7���:1��z5�]O�͵�t�����x`T^������ �^��G���$��R4�M{� /U�����ܼ�0l�ޛ�#�A�ۜx/�y��������_z�_
������M����b#����C��n�9MH�қ��s�(<�$M^R��/<�\z��o�SǏ���m�	���߾���v�?t0�ٳϼD�Z��Y' ݳ"��u�W^~!��ܳi��Y���bH^p�fƲ�v��g6���ڕfg�T���t.��75�^Y:/~ys�Q�4g��ޗ���ɸ��d���tp������O�^xN�H��-�E���L����Y�t�_ `ʪm���C~idd�������:;���Km,���Z�ga|����Q1,I*"H�%�K����g���89� �N���7���˰x����m��O^�(C�b�F�� Ęy�:��
���-|cI��XYU8���e�uu�����`l���O����Ĳ�;���Q�G��2���5D�w��wGT7w)��Bǥ0�<.v�� ];�&U��A^�lɆج�����##�t�Q���a`�1���^{��ґ�}�C�e���Y�[�8W�Ļ�ժ����ұ���΍�űl�#ȉ��[޺��x.�WY�}7��k��K,؂�N��i��!`�X#�αUb�lKë�:/�m�!/l����O��̮ի�u{.�W��	�k_�A�����`9G���0y},o�o�Nm}��omy�f���J�Ge���(և]&�M
�Ƕ#����tB�F]4l�Đ��w\�a10�{�y:�����F��몍#����N c�ónVW�{7坬�+=h��t������A&S�G>�YF���q+��L�u��WΧQy��	����!n+���,��.�����fx���$U0>�lΆ����0O�j�a4Tq��,aK�o	-(Ή� ���J���U�l�%�X%o�8�Yg�*ob�&^װ�˻ו��0x��Bz4��5��L<iÁf�-)��^������R�lQ|�o�����>06k����ӣ�.!���MLo����x&4�FR!��G��Fψ���Y@�^�H�t0�C���*�w����+�dE��Ͼ�.ީ���`����D�z�̫���a\�M�tF'���TW�bۊ�%���u�5�ؖ��쾦�ӡ�hy����\c|��L�B�K��0HG�:X&�1$����ļ�lR
��;���W��r�)�ճ���ƺ��<�Ϭl��D��3���1�]�(h9=@Y���0�8@}>k�%�w�M1D�L��B��JX3ӭu��7���S�1,uʈA��ĸy�s��Oi�#7�:�`�kJ7��yAA�bDaF%�l�Plrg��9H���My=��Pxՠ+�k�0��axm5�k������RA�x~�R�).8�ݾ�������!$j5��m�#��}c(�	�fM�R ��G2�jL�>ܡ8f{����!��cQLgy-M @�L��� KI�u�G�<�S��a�saJ����[���v8�%!�`O�1�7����@I�N��)K���ꏷ40�b)��xHx��h���e���G ����o�,���J����Q�B�����}�@�l-f|�&:+ț��[�i@�r�H��5̫�5�U��I�Q�z��g�#�Q<� F(�4�%��1��f��j*ySTA��8�e��Y��)�L�|?�^f���8�7FP'��@��c�%����%�:%K��G*� �`و&B��&�y̒#/��U���p�I�+m��yC�k`cR��P��X��W�B�ht�y���8�,��<C��O�p�3ibBǩ�ĳ(�M�?��W��d�͌٨kO浱
߹����m�:����(��<���,÷Hl�L<�9Ő��i��\�����_Q�D���`Җ���P\�"18�,,���!jL,��
��ձ d��3�k1U�m)�*��A6�]zM����@��Y����x^}����*OY��93���9�ߐAVu�۪��&Ƨ��Ht� ������0�2��=�2�o��j{���3���湳�|T�[dYL��Â�@zC���T�A�uC%���4bO��]��ԓu<Ot�����B��X'Q]<!gu��[k�W�U,�ʖT?hz�Y[+�6J���#Z��5�������|n����3��t��@#���K5���z����ц��?��F阬���r���sijvO���L�J�LS3�Ҿ��5�_���?(Τi��v�@ޓ0<ll*p֐��'�k�����E��Q_�i��(ՋgAx�I�0�s5���h}���z��g�WkH�rE�q�a���a �B�>�3���4V�rݣ�j��@�W�L��m3��{`�jO��>Ft:Xc�@{EӼ�=R1��S{bMu�IRt\nb��o��0̪����#��3b�<j���NJ)�4��C�1y.F���xnZ���p�~B��4[���zR_Y;���v��U��/����]J���8fm,G0KjJ��?D�6Ӈ0<�(�h֬P@:n�z�p��klX��"�5	��0<��ȫi_y�E���CwTJ��{yk�F�|��7�뮻�h7Z�[�q@��a����N�L�N��١��� �;Z�1X�q�c��}i��}�p5ȼ6��q#���y�9q"��,�����I�x�����T���,��J�6�|/�o��3U�O�8�IǪ�В�I�L&�$���u2���W��}IG�q�/��'�5a�ǢРc2A�B�'v��[ss���\�w��)��m_��q��D�.6e\.T�isؾ/��32���?��^ B���xV�Co���Zסw x���v`�</��f�2(=���0:��H1Rt���Y���h�}�p��+�)�7�2����cyܟ�����E�hʒ1#l�Q��-�jU��d�~����u��f�	�8��o1��g�+3�o�g�S���d��=ax���e��E8���*�9p��0�Hc������ ����2�w-�����n����a���J�"�i�^}+��*lr��Q�X���3�C3�������
�'r�~���#�ȇ�D��.p	܃�m9"@�& ��k��2=�k�c}��)�� �yt^P:G<%^ή���6����ЀS�dXf �gF$:����'U��[��آ�:������Ɔ�drA�ȀO�[[um�~�Ui2G��`�UQ�� ��g|kU2m�6Ӊo�4 #�.�b{vI��:f������m��g�g�~jff7�7Ԯ���%AO��E��Pգ���=?�lB�=uL"�ًB��l(qrݼ�b�I�C�M5��G�(��g#1���T�ZkG�� ��B	�":(��# .�\V.c &u�� W�{�� 4�f/_�ۥ8f��ԭ�5S/B\İ� �`=ۚ�<|�K ۥL�xE��xL�m=��B�����M�5�^�.���LHF�7&B�,;<��_rVe�Mۡ�<���)��D�̣z=��<:v�����h�Gɫ##J,���#N�v0Tf�RLc��s�ȑ����Y)����(�p���m�D04�BF�2�'gBs�3,0���J${ =C��pK�(o��K#0O܆��Wf�pʰ^��D����J��ϕ�9�1X�s�\�m�s��j(>PFe\���R9h'��Q`�i���+�j�b��O�#Oې�+��ݒ�u
��DId��x�᲍���u��h�)ş& �(:���E���3����@�E��r!s>ˊ�p/�3nC�!V�.! I�ڦj͉�ͷ.<0ܪ��&�#�F�Y(V��j�
��N ��bQ6�1�͊��Sk<�3����|���#W2�#M�FԴ;j���V��G�< �@�aL�A'�W��b߾��`��&���C~w�P
m�ǦO�:A�G�1$�O�J9�,k���TYK�%@��̈��2d!3�E,�x�o�-�m|	�%i�C&+k�y�2*�2^GP���F6�"�~[D+C�:��钺i� Җ@�#U�d^���a����
`O ���9�林 ���q��p�<�<w�vw ���(���͡,����G�{~tm�7�2"����F��H��и3z��a��C$-��+�$���"kb>y4�p����U�m�pr޹�/���>R��/���H�����0H�_�sJчu kB���dd��
�b�e�������z$GU�?��ŷ̓nx����_.�d.t������S݈��`���`0	ӽ����-���� ��Q���.��x�k0Z��x?��r�v4�|��ឺ��J���3`J�rx^�o{^C�6��q�=*i�9^�%/��C"���\&��h`<���|0Dk�གྷ�r��K_�}����e̠ttC⎇�>�`�T}[Pi��3�A�X����+��@55�LGO �b��>�x?C]�}u Jso���R�Q��9[� ��,�i��9^a1�y`���5DҸ�.ch�&Y�R�;
�w�2ecf�Ǳ�~��?�a��+�YRRl%��i�e�*W۲=��|�����0�~G`&C���[9�!�	ys������1��F?1�0�xe<�����1�:_�CZ�DE��rY:m	��y������OCB�Ƌ�Qi6�w���$�f5P��YSuʳ	Ɯwi@�#�⺚��/�[�j���P����;�	��׆AKik�8�]��Ax;�x���Ҋy0��L`�W�sQ��H�B�� C�KE(�A��?�,�-�z�����w�qP��	��u�$���4�t��2�/<��gu��h��hx[X�5ʹa�	Nx?�#�鼞�6�Fl�BG �1cT^ҭ��,�����&vN����c�OOO������gum�2� Y�.	���z�
@���C�1
�R*� i�@��vtYz���Kv|�1H�R�NQ0�͸��f.2ІZgoǎa�H�������C%�R1%+���pX�{���<r0�gmb�_�f�feSAG����M����	y(�!�n�c��a��)H�h���˳�,YK�l�`m�c��g��m]�^d<`D��r�O���E紑=zx�QM�x��0dD�Q�UƘ$yxbq����;��E�.A����Q?F,9"D�eCBf�	�;�������*�<�.`�y^��LEl@9� p����pȇ�cϝ�����z��Y7x�1Z�RO���k��5aI��Db����E���%3g<S�屖�{��ݥ�,v�`~�FhF�Ze�t�s����p
�vӤy$< Kt�<�f���?"�#Q��H�e���"�O$|���@L�0��C yMb�g��s���&Q�oW���Y���u���o�i$�'��%��<3i�K���7�����듓�_޼�#c|��x����?Vϻ��΂�l�����t��q�� &�'���1x�x���l�rg����������Χ����9S(a�uz5Z-�򇠻�����_�z������oM�oX�c�peu=<|(�p�M��2>b���+�S�����*��W^�����.��׸U�,�����L7�xK���5	���K)���>=�Mi�m\Y:g�1�.�Ĝ�㣶a���bdo��_����g���.�5�m޴m�>}��k/�g��uD.�L����V���G��Hk��s�e�1�Ƚ\>���96�CE���������	����;��v	�cb�}�j�d|w��C(��Z}�nW�={&?��=lB���|���G�Q[��x���xvo�&��;�h{���?�n��N�>�v�0t���������'O_���imu1�NNf7�Y��:جj;E��[�+��w��]��+vlxL����nF'#`X^_]N�<�@�����w��NN/X]�0�#�z{�L�~�{ӝw�-�KQ�dI�b?s���ڒ�w�}_N�>���W���J�oR��$������;�;]w�MR��&�����M<�[x����/�g�}*�<~\C�3���l�Ok�w�o�����9��ٽ�R��ە���o��Y{o�mN�"��v���}{�۱�������`����0	S��U{4����S���3K#.Ȍ�D\�؉�h(ܗ�ʲb���l��9�b���:�+eCn�UҴ�,/���'O��G����_I�����?�Ο:�E��=����O������T�x���+˫iii����x����si}y-����'��˝L���&�A��1cC���%C�)�zCr��pΊɂ�אoU�0� -�;���8�ݰuٞ�[YZ�n��9�7a�㥱�����^V}�T�R�^�/��OK�Υ��E�l�k��/O���T�o+��ʊ������3u3��!a�s�C�T���%�s��s{XE=�^5!E#|vI�Ƣ�<(5����DJ��6)g��ud [0��R'`
Ξ+�.�<.�0\�+H)P	��0����1d3FІi��ҙ���Q�:��)^q����ϭ&��8g�Eg�`�!ed@����'Q2PՁ��!���#å���$L��U2�4Jț�{ß:�r�Պ��Sy�V�:���'nj;3f�E�dω4�l�Y�dn���E&?`��N"������\�Q�q��v��<��Q�ժ��p��x��0cP���U).�j�M;�8�}x��M�<H��Ca U#d�]Ð�}�t�e)G2`���A�x�2k����oGm8#��o� !Ȯb{�����^^ZW|+OU�62���S��S2�5�d|���\�Q��{�P����#�ۋ��"H���2Pbc�0*}���+*�9Co�'�ե� �B�8��ݿ�Qs���w	�A�Bg`�چ��`�o��Fj�EW�l��M�C�0Ƨ G���"Pr��1C%�����ah���3]=��t�=g5���u�K1�@�y��]�G6�Ѝ��a�F2\�v�U�5����.q*���D��-<��[�Μuӯjx=v�dz����O>�^|�e��11�,�(734x�i ����0��aϐ�7�'�PL{9�yj	�:���,�1�Y�	�9��҇N���3�� ����5��gT�W����Si�a��3����,ίm�^G���Q|jXKe�+j|,2O����4�����:� ���1��T�b��Pex��o��x�!�#w@��%k�e���T}�$uK��=ou	�<�`l��e�|7留/7�)�oN�$C��.i�I&U�m�W^>��NA��/�'�|6���񴸴fm��������Q��I�x5��"�:�U�T�Jxm��#��-,ä��ӌp�D��P!�[�q����;�{M�藪����Sb��o6�v���;�5�9w��S.�G]�h|kkke	iB���c"(�a2>�Ȅ(��Pt�f����76���Q6i�A{LFų|���c�s�MMOe�>r1��x��h:v���iT?tm?���)C�K���fM<��:�_��f{&4������� �3��fI���%y��t�̹t��U;�_Z���y^�,��Q+mn�,V��©c�$y�v)-�)=����d)y�ۭ
���gy��ŧ��~K�����Fm�p0΢:QIm���
teZ�H�:2����G~V�h��D������t@�tŨ�0�h|��N�3��Wt4U7�qC��~ۄ_�B�,�FeL�vq$5$�������%�T�P��dqTF)��H��ʸ�N��?#J�`狀�u��S��L�=|�kzm�����,��O�I�}5=��IO�5\�r�tZ]��Z�ød!�����0"�WH=�PR"�?�!�<c�_A��Ԯ���u��ApS1�)n�E�n�P�|;��v(��k�6�	Xv��T�"�K.��b�O�Mȫӱ���6Ĩ�DV�{�;��-��{�[�����Q�n�� �>�Q��v�$c
bl�@'d��rxL�.Kw�MG�⩶v�Ɐ��P��ۇl�F��׌�k��а��ɢ%���m���������vV�q��Da�(e��@],ңg�H1T��%4�F�c��*J�fdL ���N��G�L08��VG��H����{_�b�엾��}����I�>�lz���3Ͼ���8��W��1I����^WA��(o�2���L���cxg6}����ʪ���A*N8 ������B3:񎧥N����, �{9�/FF��h
�j��|�g�y�C",��1<��1&�]-6����t$�S����6��	�;�e�E�>h;�Cȟ�/��eB4
v4��zf|�cO�ch����'��b`���4��x��φ��	�EU�5Q�i����i��C��kӮ�=iff�3y�-jkA��8�_S��P�W�{�x��'�lqI���45=��&T�f�#i��Q���B
5��8T�u�G�Ey����[o}S�����#���#��5�Ӟ={Ҿ��R||��<�f�Qv�S»Ő效�eg�<���8�����">mK�dƤ	KC�bJ�V]a�8�g���_�d�Cy�w�O��.�s�܍,D	=��ّ3�c����)��e��-t ȸ$lllhTr����7��#4΍�!5��J�\W˰GR �0�����L��c��P9���̰��x��T�y����V¹s����܁�^���Q��a�����Ӯ��yl�: �C����ˋ��ٳ��i����7���w�������~Q6K ��x��.{���J���Mf�K�e�*��6�	rrzƌ�NO}�.��ʂ�&&���K�Ο5C�Y��6(p�����'~#;�)kz���c86bG<��؄�w����`߾CA���� C_�����j�o�G`��$��6��rB` �s{���F��g3-����h
�::y����z]I�v���>+S9�ŋ0k�df�����%+�thF[u8m���gXa��Yb �)B��^�F7߹�d�w2a���X��8S���+i(��䐎���:[̕⩃|����aTm1��Pr �09��M������7��O�Ɠ���䜴�!��yoCH�e�.-��	%m�3�߯���G��U�+c|�E�ۍ��h6?��6�q��c�F@��L���;*�0-Α����V
��a 䥡��a$fS͖���Ŏ��>l����"�X��.��6�"#���]��6:���乆QX{�,nWYG2�ݻ���#��4��+�;'"h�e����ר�|aZO�,vu�����*�FG�#�����v~��܃�@旆c��^}�t1������ۀkj`���0 ���V��X�f��2�-G���d@G0�͈�`E4���a�oKfD�0eV(B�z;�u$F���C/��ڋn�����(g�{1:�6��d�=�ģ��q�hRw����"d�� �c-u�`�&2��1�&�uI�k �9�D�� A���r��?���_��{JF8.s^�u�N�@\�2�m�?xD{%����o"�쾩�64�ŝ@�'�����W,�� tn�lU���Gǰd��gH��@y���q�a���]���0�V ���m'���u���#~1�'��<Ц�xC</)��#	�����@�ϯjc�K��#^۷8�'-��"29�0�/Hg��A����cD`x�;����醎Al�f��
��,��>��S���'��<�\3�S��%;��L�:�Ƃ�p F��j��] ��<����g���ƲrT���%?3-,�Z�#~�=$�6,�dC�����o6�L�yF����i�]1�<f��Ɋ3�4�cU�w2kevͻ��	l<�����Ȭ�0PF$b9�o�%?#��3��9�v��64�Ptt�Q�,ˀ�axc3X5)deE$g{�3���I��1�m�������s��h�џ���?�����R�(���ѣ�x�@�$b5fU������ ��(�Y(���(D�t�]��D~~G:6��D�_|ڶnd$BL�/�;����زE�����Q?�`#~C%�o
�ʲ�2�ƃ�$`��Ob�|���H<>��ϫ۠�lz�)ݔ���s�p�g Zf��v���!�V,��Ay�u�4�g�w�$_]�������D?��F�b[��D#{��uf��][�MhC���Q�u�kܘ�<�Qy���>��ǈDTh7�u�T�uz���7å���>�x"�R��-a@�m]���Ķ*޹�anṡ�1�5�cA�B���y�K�*�r243���aQ�w s�<�gO驍�?�[S� z������F�;{t�؎���E�� H�00D������R�ԛU�H�'"�xn�(R��(0J�E˞�E�y���ƀ�n5rx����+�Ut�C���#Je�#A%�D��𲖊a�����WBP4��B�CÆ�)L���<}/dk\�̠ ��2>���'��$��tD�y:��ɗ�٭��P(�4=��#F36Ƃ4� D]9�<��S�g��F�ol��Y����0x�eh��V�huX��@C��ϼ�Σ�ὁ�;��\���z%�FP�Q'�����OeF��]j���l�K����t�v�̩'���-߷�`ǌ���j�'[��ߔ㹉�h���#<���A�L8ʦX<�y
���5��<� y|��m۵�#A��Ɍ��V
���m�3���E�S:X� 0�"��� ���*�"h?�NZ�fe�����h�s��#7��b��=����^[�>���(`��Lx�o^��Fe�D� 	��h��!�C}�2�ǚ�&��
����:l)H��:!��Nd�*Fo�o�v㫳s����}L׶�ڋ���N�m�_����X��L�55Dޏ�̓��(����3�AD��t��q>��F�G�9HG�(�炒�0! X�[�:*,�(p�q���xv�vfhx�ժV.�b�R��	&�'�C�VCe�׬�.>��rj+i���09�VWΧյ���bxd�9�Y����w��C6lk��8d��itj�����x!7�0*h��s��./u4�g��ʲ�*c*#���#��������&t������ő�L{*�+�+��Iy��R�k4������4��R&�B��|��s4#���� �Uf��Qw"ڍ9�. �[C(��[� r��Y�ńx޶��q�WΙ!����J@�7�ʹw�>{��6�k&+��������R1:QqF����� Xa����:[�}I�f��۔��P��n�j^1��|�m�,�Q��x��꧃j��2	���-4�H��LI�� ����Y��zvM��n�CuP/�6��\�� ��9rQ<}qzf��[z{�2;����1��zu�'۝��n��}R>����6�d����_T�i�����h*ckI�b�%6�n����˦5�"�Ç��W�<xH���Ā���ڕb�K/���q�yqL��䧬ߋ���e��ֻߞ��ֻ�®=&KR��"L5�����3O�g�yFrX��:���'�]Y]M�>��:�D��?�_��n�S���	,�@E�\2�Ϟ��fzⱇ�+��dO�q��]^^�{�<�<�#G�m��fr	d�e�j����"m����t��r��
�>�g�ʑ�ۃ��aY�,�n`e�ƌ��+����<]ȑ�]ҋ��߆�B��la~a�_��=C�����O�~RF�74��dO���!�"�yƓk<2y��Q5|�i=���Ĕ��%ዋ+���kdl����ϥ�{6;��=ų���~w��-w����m�n�{�
do�
�C�2>���7H_�ʗelKJ�cq��k��@�|V�g,�����~��i��k���h�
�PX�!%��|�K�o�'����$py[>-e�f�d�������W��}���?����{ޙF�&�[�P"�1�����gL�_���׿~��(F��ϟOG_~)--/��p�c1�=�yO����:�#ڼ����)cS��c�1�����:}<=���2�Ӿ
�-Eџ����W���E��t|��06~�l5iȚ2{��M�2>td8�ٸF4��Rm9�/��G�Y��
��L�;N���=���?;��� �6#�P�%�ɴ��9	��t�_I_����W��8ހ�V|�!�M�T��.�PˠT�5\�ӫG��z4=��c�O���~:=���:>k�����'=���eY��A��c���1�5͉�'�/� ��h�	�R}/ۣ��w�yGz�]w��Y�#v���O��<%]G�A� ������C=�����ܳ��3-<��W�ϝ=c�/Z|��F�.��=�&c��x��j/k��T<�be�}�����pi�d_]^R�Ey�9��P���yΆ6�5{��cL��J��j=xh�����)D��r�.��_w��fA�H��1���)���~����7��M�gҍ7ޘ�򖷤[n�ņ�]�vK9�g���,Ɛ -腲~�~F8ƶw�o��������3�O=#c{F��S2�^�4Ο{�����T�a=f�{�Ař���./}���ǟLO>������貍kc�?�޾�{��
�Q�f�\@xƈ-��|X��ˎU��3[2��}����h���<}�#���':t�<ƆLQ���I�!���J��x���nR�p�g��7x�t�i���u0Q�#��i���B�uH���䌘涽7g����j�b*���Ww��#<��c��L�ꑇI�+��%X��x+��<����Ӷ�ݔ�l�f���H!��j:{n9�)�_��F�Fڨ�<�<��0Yeȅb<�婍��>�0�뼼����^Q�j;�	��z8}��(���4[��Z(�� ��۾����	֡#��7�hG�8�]�yw�����Y�ff�OR@����4�����-�����k�MW�W�7ʂ�����vxM	�dK"�š`G�t��fQ�f0�D��j�f�~M"�p�,���������������O�'}"=�У�%y�եe{��6`��ԅ �C@���v%�a�sf^�uXĪ`A���ً��&���M��PP�.��R��]>�껇�h&J�;M��Ʒ��?Ȥ�N�~��{W-/ޛ{�F����m�K�v�aN�@��C而>�Ϥ���Ӄ?da	����D�e ���'i٨@M:���7����2�����M�|/��R��<��)�~��?w[�@q �;�Wr����~�0������fF6d�7�,*3ԓ��^z�e�D]�ǎ3��`\ �а������0�0H��@)o/�\F�bx&{҆#�ʃ I'��Cq�x<��~C� ���m���1pv�2��<tuD�����-t�;�U�fx|ꟻ<�Nl|�������Y�J�z��IylMH��ųVI����T�yn �����nȱPn!w[&B&��� ��Q굾�5��_K2C3��!�gTI���J�"���w���4!�@5<t-��zU�3��� �" G��xcQ��943@z-�F��>Ȭ
���M����'A���UŅ�'�oru��-���MIY��}~ą�E�0��B�B%��,��m�uڱ!�odE0��,�}���Vh30J�*KS3ӽ-]��x���'x�_7 �Mu���C�2��>>� ]��f���D^�Qdב��}2��`�7�%^،�P(:��cO=���+����x*���5d(��'�4��n�N���Um���ĉ�&Xh���"Yz`
M�����` ~g�u!�1r�͢�hI� P��(KpaȠ=�n����糸leT6�?S3�i[�c���6ۨ*�1O(I���^��A3���ch���vYlT�f�I�x\ޚ����������H@L�+�F�؞>y�B�L~�w7,{[xE��s���8E�'^�t�-(�D��!a(K�v[�p����ܨ������w�!hx�n��|OIyK�f$\vIp�xG׹7�{�v)�ޯ�����&5�1"�W����̮�߅7-�eD���)�˔k�MM8�W�Ӻ���$#_�Lk���5�������ݨYB�C,..�^�6xbn#�W[�(� 3h� ��aɌ��"1"��o����;�3��Eϝ_��j�ˈ��&�y��Y���21�j�h����x~�l:�`/��C�
��� j��G�p��xD<��UX��n^�@�|[v��cs+��M�x�d�喟pl��&[��6 %�ml�~hc���f�-T��j1�7%t��4�@~+��=GC^��4����'N����4>:�}&����:�b���l!vaa!>|؎���y���~R����z�['�����S�Ed0(c�<O���}�E[���d���O�[�����~���_�BZ:�����)׈e������b�G���>&��'�z!��Gf�\����^=s*��o�fz��MA�n�bV�N{�7�;�+]{�w���Ptl2�3r� ϼz�^:y�����[6` ?�P�L���f���#_�q(��"7m�!Xh��i3�Xa4�}SSӵ�ɉ�޻���Gy�g��1�))���Z��[���[�}�1E����PB�G���S.�@�����у&&x�LC�z�Gc@��!�LC��P2�L�܈��0��iD�����c�O�8Ƴh�x�چs�����@�zϞ3�_�*B�Ȣ�Ч�Dì���/�W�x>�e��3�~���_��6ʠ���tb�p#��dw���1��}&�^�Ͼx���ЌV6q��m��-�ބ/No��6�Hh�L&}GR�: ~�3��h}|b�Ӈ\����_4"C�0�7]�o~`s���N�}�*�2`�Wx1�gaFX�@�&��1��!H�kht����
��`XT�T���@?Bm)Ȍ�@ �B`����� �8`�U�-#�΋+4.e��x���8�vK��0xd�kb��x���ƈ�ؤ�ڬ�Q�rtf��Z^&����(2�<y��q�9�!�{�λ�)Ϛ,�q��V_�&�KY.��z&ӁBcll�w�9r�
�X�!�_�E@�O˫|�^�~J�߭Jꕡ'�`��OƼ��t�W�!��`|Dç	S�LM�����hl!��&;�Pԃmc(�$(��7 f����O�.� �f�H��YQԅ����ɤqn��
"/@�e�6`�%S&���S�2lq2O��8�7]&!�����[t�T:�ڒ]#����2Vu2�G@�~[>%�������P�Ȯ���7�� Q�d�����U��?�0���e�Co,p)^���,�"EL����:C���b8o��-��
4�Kcz�tN0~44`T�QI���$��F1�ztF�1�=C�~�s�k���B� �_ĥ ��wl�0�A���oW(�#���N���l�Z#G�͎�Ηr�W<^ ���@+腱`N�҉�:�yM�ۃ��Jz�>ґ��@6,����T���¯ɡR)�ȫ`� w�a�O`��.Cy ���(���"h��Ęf��(BG)�5�#Õ���of&,�5!��cuPw�_�CG� m(P�"���j��G��=�M]2Z������?!!�����x���,�H�
��1p � fP*ƍ�����QJ���QG���z�ǓifnF;x�|ɇ11+4�S9&�x�0{&&�)���= ��)o+*�t�,ޏON��:m���@
����P�@����Ԃzh[�%��!0�� ^$��Z�q��L�1�1<ҸrNl���\z���1��)��tĶ-���U��G��/�\h�L�z=<`���"�6၆W{��a|��諌�+/HG�ˣk5�7�@�<����c��4����@�����h;�uB����'cdb������%=r���X���t Ɂ��xFd�%�1gdHت�@�4�)ʓ�YxH����E�0��,H,x���Q�5
e���VA�9�RɈ�5C�a"�IN��))�QPG(����0i��!!a��J�)�z�֏�Q��gó���S��~Ǿ2C�x+0��<���c�"�Y�z���S�E���$� � �@�=%B/�̣2q**�H�0�<��x�h8���$/�}�eS[�R��pk�_��.��,/[�-�t
���%%���V*8��-̲}E>vg�:4��@�ײ{�	���Kn:G�ރ�611�B�A!<Ι 0��|��ߐ���\A�:< i� HG��Ȇf ��^�<`���h������ybxI� �;�^�T0��"/i1&�2~�t<�F~�\E������ǆ2`�m�H������D�*j�\チ���:2�a:.�z@�WU���)B�R���(����Q�U��.�!�/�K��N�A��e��vgJ���z��B��#lC�j2�z7=�gZ���k��`Ix|�
d��xh�7ҕ�o�?�[��d�|_lbl4M�|&F�R2���B� 踏�k�#�fԼ��/h��DN�B)�3ɺnϼJ��s-�~�B=��M��7��2E�K�A�Lů�u��h3�A��.(��VE��I�O_�	�r�^$3��;������3�����Gx��<�\�,l�1��w�1�!A�/j��;�]~Qܥ�t������m�"gZZCq\��4�����W�F{�C� �7���dÕ��Wx9�H���du�1n�Q�����2^�:"f3�e06)�(�-���0z���1�$�٧m����0��dб3��4����l�,q�	_��iFxy��9+#� l�e�ɚխ����è�*bG��C�y�6Rp�sB o��pJy���<�{�OE֮���f����Wg����=e�C�s���J����
�)A�eG�YA�&E�z���!�t�g�5� �����1T���S��U�ʭU4�Fz�)φ���-�.È�C1���Ĥ��@1��2&&&��^�'qK@=��ש�x(\5��dO�wR~œ
������3�e0(��&�y]��е��b�"���a3�</�������^1�:��� �)�'���GՒ��}Х͎����WW��7C�U@h��S��0h��=�w�I��^����%A�V ��F���%��L��x�&_�A@B>Ӵ��l���K��F�j���X�#���]��⸅�=��_�#�R�˫GK���~)O��!�h	C�@�e^Sr��+��?x8�ݿO�^4DWYz���r��.�M{0�� 0,m�،�R�xb����l���i~�n��`l�������K���x6�^@y�|s�PD���\:x��γ}��ċ\�y�L��D<w��6�G���0Y��l���s<��1�?�kC����	��Zc�\)�������h�j����14[�V?Z�m��ιá!��@���"a������	��9����`Ua�EH��Fz�]1�q5i�ظ.��K�[ޜ�g�L��BH�PYy>K��3Ϥ���jZ<N���I�E�m�<�V��lm�'�n��N{���R��3z:S�3"�E���3O>�Xz� .@ѿ�gҦ:�$����� 6N�,���Lzǻޝny�>��K2(1{{E[r���+�_�|z��G��ںm�Bv�>16f� k���tcz�{ߟn��Q�L]�3ؗ�$G��x���ӧ�q�Eu<��|��o|�ɄiA�d�6�S������`�.9�` dI��-�)C�|Ϗ��������/��X%C��Ʒ���V���8���f|<ը���s���'O�Fm�&4Ζ�^3BP�<3 	������W���ѱ	�;Ҽ�q�V�3:��R���H��}_K������	� y���\���{���}�xz�?��g����T}����������/�o>�@Z_Y��0��W����ciueM�iW��� ���԰,�5f�~��یҹߊA.--�����J_��ӹ3gM���%Ϥ�s�6���O~��o}�չ���cTʷM�xe�#�,�ҋ/<�}��t��I�(0A����_��~4O�7<�׊�a�a�ey�i���yA���O������NNL��{�L���1>���$� k[��(�#=��������=��x�!����������m�����.�U�|f��ɪ�~3��9z������c/�x4�z�d:u�x:y�X:w���{:�=`h�X�@a�8]�p��S�/c���2[ǬY��o�*�<��<�v(�4�.�D�1��6m'?n�1L��F6�z�8���O:���)3oEyx��aT���) �^�PO�"T�TH�!/�����{��<�f��+��rN�=�r��������0Lf�
:s#�cyâ*���2�X��G�)�#a&�a��&�rЪɳR�k@G@�n����T�`RC �P�ьkb��;A�������4�#��	�f�A��9�G��-`՚+\Y�7,)v�]�ɪ�m6ÔZ <���N;� �s
2`tt��ŀ[t�D<G]�`o��[t����nב������'��ɝ�L��	 9�<�P26�⋉iy(tJP�ˀ!-�[hK,�0����û�^��@�mk�0�4�$��O��0 ��B�3����P��5���7[\t�C���C�&��v���� +���M�0���3�za�/=�3�WQT�7Ҋ�{��F��y*om�� �Q�I'�Bş�L���⟙)3Td�z�T_�\\���...�S/�?Ǒ�e|
oD��#��%λ�O���M�)�P���m�NY�gR��pD�F^�Y��1#A?��X�n<d&㛺��g5�,^��qC��Ø�*Ë�{�vֻ#� F��7f���7+r���{�D��	��M���if��N��-������Ef���K�4SEN�^���!^m�Y�����U?��;F��1�rɰG(�k-L9�:�X��l˩��KG.(T8��=@�S}��C�����!K�F�O/�� �Q7�`�Icv�wC���­9��ֹ-�(�r����G��N���-2g	���N8��"���^n^��	9A��<��f�,���[�x&�v����Qn�s���x�B+�F�u��_o���}����p��tN�O��P�A��(.����,�����xxhlt*M����־�$o:/�G5�.��r�f|f4H�zQ�%�(����?�_K�k�iM�����D�_f����9��Æ�dX[��ވ"onw%�������ɨ?����!�KQ������aK���˃b�����8t�[�0� �Z���nK=A S��f����G������<Z�k($v14����Q����X]�.p�!�M�,�x���AL���N���i�.��[{۵˟!?ʩ[��� �ę)R�ꊋ��L�mcx��q���}���,�G����
a�Ҟ���=�D�[ޚ�ʰ�k���5y	�`UY����Gd�u�ѓ�h��gwpXȖ5��]�S|��Lo�m�2}���ЙǕ��q߾�O_��ZY�)� �P�2H�	R����1$b���E��W���zy��4ȓ���b����z�"P��75$I�<�651���S�$�ci� 0p�1Āh����6��q�����"�Y���;\�شj���[�-?�:bƿ���n<��4v��H�&Zd��#��d	�ظ�¶|щ�QY&aT2T��
2!?�x�F�&�ڨJz�!@hM@�];������:P�m��-.�!a(�W*���_u��ְ��Qo�+`1 {(Z9A�3D���Q�Ex��̴�Ҭpr&����;Jxw����Æ�Q 87@W*�ak�i�����c˾�R����'�N�|��FՂ}��o �Rq&
i�WJ�J��[�M�^<�X�����(�A�(yP��2�0�'�g�7�GC�3��Ec��Y��)ތ����*�[t0Pbh��<5y���k�9�Fw�"�͆���ɒmf]�k���^��+�s�F���Nuzٴu>���!/��2۾8�a���{�7�Q��۹���m�h���x�	K�
i0~�+�")<BB���Bz�]�9Z��8������.�g�Q�[/0S�0����^~��t��R kf�by v2#@��CG���o`�T<��5o��#k]O<�p:�ҋ��_�iwN$u:��o|���7�9�x�-��,��o��£0{&�W�6c�������/���C�'!?�d8��S����}(]����,L�2�p �{���ԉ���C����=j��rK2�<wf@f���I1��-�Pw��T�����O���u����{��ޅ�.ھ(9e|���{67k���4�@(,?��?n�[���P�:�Ćkd�e�͢x%C.��D�eC�[��7Rr�A1[c��p�����,N:��@b.�,	xH{��=�Xpzjք�Q2��@���͗���-//���=i���cU)�'��eLh�1%���r��1S�]����B-��C^Ή�8'/�I���-fU�M~B<9�+�nv-���1k�,�[gґƓ�B��5l�y�h�GQ�>��V$�ٛ�����F���>��k��ٻ�Я��5�I1!���Ey�ۍQy�]	���}U72�S�1�3��#���L0�Ȱ@9�.��1aI�P������a��2�׃��G�P(#�:Ʈ]���(�oz�긥���y+�@���g��w��C�x�Y��~Q��=�L>r-�Yxu ��uv�@�� �r�6�Gk7�C�'D��@G��^�W"5?N@^гgH�Y�)�0�T�8S���3s�?#χ�]�z��tq@E���R\,����Ŭg�01��F��#	Xj�=u�{H8ڛ����5�n^�oG�@Ң<DG�PPjO���x+��*^���X�`8G���'kC��/؇h'q�ؘ���7��S��	ĄŬ�ɀ��Ex������aA�d(㈂�!��S:2d�7<'G�����\B.��9S�ʪ�& r@'ǩZ���0d��Ѝ���J/�H���'߈���1>1����׭�Iug�ٚ��b"J �v�dȹ�� H\�;�u�=]�t��@�p�i����N�@�=��`LF�N!u�u�W����{t$�r��(Hg6l;��w4\��h_3�@�2>3�^fv.;�E���=����*Ox�Z� ms�T�*���0,����"#�
�F�g�lybм�t`�pt$��|�:���k�2ш�T!�x{̕ټ��s���y���>�ӉE��F:�lbt��[�0��)�.��޶қ�kp�^e�����y�L� � 
eM*��,I����Κ�o����#hKBf� Gfq쌡i���10h�n�/L��Gd&i"gx7�?�D{�a)�g�9d�x?<���G��O��t̃fm��kJ��F�c4A���_���KyЮïh�Z�����fKn��|�\T�ȵU��D�M�@[�6.\N��Xǵ�����/�!����ab�<o��!/��$0��a�D��=Zh�(?�>u0� �(�À54@�ms�D�m,{�5�+}�!���z8�1h�hF�?b��w%���w�h��B��#&����up,;���0��e���q�vTG�?�J�5�c�r�y��>D��(2�����ٌ�VT^\����w%�f�o�\�s��H�e����MM��Ta�iq vM���?n}�#�_4-&�B���P�!6@(�<.4�Y�9�
F�Y[EW~�`�<ই�FE���q��m��+�-Oԥsx���7�A�E� �۳���>��p=��s�y��Z��?_��͗Ц�a��|���>�T5�ݘ����&(��7 ��%h�V��K93d�����m0ʉ��� �$s��7�����9X����O�Ƃa���-I@0�@��@YbזV��VcFu����s��Y�f��h�`�w��
�u$�3�^<�F\A9v�������B��O���J���iK�~���2rYM9��]�q��^m��YҘ �S~vR��r�,C)�ZlWR���=�at6�R����g���TO�8'��.�Vϰ��c�x�"�I�w��}� �Z����[�;ȏvif\aé:Z<C��uɗ����=P�c��2_&%6� ���4H�j�ݭV���w�2M��&���0���1��������IeD~�
pA��#Hf� C�E^�"P�:�V�r�,���� 
Fev���Q	���a0^,���@�ÌP�W6f��H�����uދ�h��!��`�c-��A��8��=��c���j�������_��"��td°/\����eޟ��]&y�-�Gh�ՙ)�����0�S�Q��Tu��&]��j��ё�ߚ�����ƃ'CA&�K��!�[�_�D�<k8�[��=gdL�WM�%�U��w�3Ji�V��:^ʶ@I0�`����9'"p�����O�ؓX�Z�RԐ��j�'fI��ݢ����hMhuJA!`D'C��>�,%�)w�����4+e�*�W�0�����g����#^	����`�d�M�@�R�{�<�-���6*I�|��l;���X&�7����F�h~�>���̢A�S0umFB��*�Zzn����X��,�7��rn������T[[N�چo,e6_h���|
���t��A�=BIL� ?Ñǁyc L���b��0˳<;���Ϊ��`�����h��cu݆:�pB��g=��)d�ԣJ��y�%��W�ޤ�x�=u�)۪���j��ic�\�\]RS�n����4Cb�0�L����y}�	��o�^�[�j�#�d�2�}�cG����_�49��]�� ��c�� E�uΑ;Ft0[�U�f�eI�ޛ'$�Oa�X�c�%����.�K���ɭ�]��S2�w귂�:�p)������U�{/[���vu�;dD�ieձ1A
0��~�d����8d�����4Gi��ި��~��S�1z%���A�Z��S��溴��[)>ąa�h��:G���Ey<r��	�&#x+5P�鄶�@Ƚ��tk����e(�'^��Ŷu�B6�^{����s�=g�E<K/�=9'Tx�-��;��^� h�e�-^�������a{y&�W�953t���u�A�q@�r��|�_=c������y;�Lt{��u���c�������D#
�2>	��ju���C
-�tK��n�ѓ�}�������	�G�Yh$�j\,���6��8HQJc�`����=�;ߚ��X����f�B�3Ďi諭���y8=��#V7÷Ŝ2��c늊�� ��oW��ƛ�l����9G������}���?=��#��5"��h����(�����g�����~_���|�I���[�ˡ0{fB$*R;���/���{���mxų��#���i�'>���g��M7�t�Y>[�PݰM�^�#x��'��=�N��ëw&&}�%J~҉�ˌ�]ጿ����~;_��C7|�/F�_��ܙa�̤����c�SS?93���W���k��{j���7�{��j�^�-��i(bx�\�H'OO/���y?bG�+�nt�`[��1� X�[p7�Б��?���{����I:�˖�e)PIS�%3���_�ڽ���@ ���]e�|l��[���J��G��w�m�Ψ��I�N �s���U�n���?����7�~�{Uu��h�/���wh�;tM�c�ӛo�KJ�Ұ�0��ty%<[3n>��O����>���M�N��z�|�cBC������O���W�J���[3���3P�@:2�8���=��7ӗ���t��q�i}�T�leA�y.Y�����2�'Lt�[� ''����]w}���N2<�d}�����������ss�O|�n�!��a�P�`��Ĭ���=C�Bm�e�eT2���\*V���Elё7�G���b^{�CQ��uq3`z�0$��8J	2��-�4�lSq�����+"ڊ]��A/����' h���Bx��e���b#&O��R}X.mw/���L�ԧ���N�g�w�J�Ksx&i�A<�N�k��^$����Xax�m�ZGF��SgĠ�ȧ�-ɕs^�n�����i�����|�U�L�چ��'Q@U˷΅�P�'^_vvfy��0�b��?0� T���� K����-����#$�#��ϻ�XZnx�����+��Ф�/cC�@��-�g��'ߩ YQ��8���A2�2�`Px�fmC�4�F(��t>���n��;�P���Sb$$��#��TF�[�(�'
�>q�dA�����Wx��kd�p�����f90�R;E�Ϛ��M��{�Ӿ}��#�Ӯ��4�^33���9��+��d��t��k �<�K,[�����|Ϙ���]2��:0#����:#�,��ES����[:�76�j"��(��:���:J%b��a(�k��n�]��Xϲ	�BC�=�/e�DC@,�3�|(
�"�����
M1��l[��*Cb��b���pP��㜅]��n�bP�=q%Za�<s�?v���C�=�Bqᕀ8'(篝+�2�v���1������)/���=β���&_������af缴h��ٴo�B:,/x�ྴ�.��M���M{�g҄� �1�X��ꉺ�.zrS>[Ȗo(�� ]z>���9Q�d��$�ͨ$����+G̨㦁H�6�l��]�9�b�h�'��hXU�f�?����(f�� ᨈ�>p��� y,�l7$![�7V׭�R@�g�*�#� F���q��Y����>.�,!����l�lt3�G�.�L�Q�%%bgK9����Y�,���4���ӕ��`�DKհ�b��S�ϙ�s�KՑ�6��޽�Ӿ={���kN�v隼�:-H<���y7H�t('�-���m2�Ei���amϼp���2ػ�u��ё���б6$ۈuy���={V��]b؅��Mf�^�8Ǜ��yopٶ%�&�2f�$���DA�2 )��"|ц}b�O䦶�-7��/��=�S���۳R�MP�H�n�341Kc��B��,����`��߆{��}*˰i��2܉wJ��(0�o��ç�x���2����[��9)�����Iu�
7ID�prΈa|+�-*	B��f��#�@����#�C3�C�Ȉ��}Y�w�R�+�4Cy���CH���>���.�0�0�N�_�i�j�fa�0<�E\D�8TO0�C��j�x���� o�����#�Ä����sBU��k�S�THؕ���-\4����vHBv���i)gܔ/�J5ʯ����2>�6�l�573J� m��:�`|n4�S|���*K�9����i[���vdD|�K�v.�Z,h�a�T�lTZ���	�;�C�	c���`Y-�����z^��Ďx'|1��n�����(A��;���B�>�Oн5_FgT�� 9����/�y��2U�:��&_Y�qc�����?)v4> ;7� �z��8�x��n�%Q�X`�c�?Ʌ��@�+m;�u�Q��Ɗ�W�v ��A�&P����xS��o��lߚ.8�B�q�"�ҩCyX��0:Fߍ��5�4t�nxU�bΰm�K�Ykt�FUʐǥ^�P�{u�.��ʍxd<�ա4:B�c#��]y�8O�ׂo����G#:'V���3KVx8��:�[m���P��F�<-g�E����9��?�s�#@.�'xu��Bv4>Eb�l(�	��߁������`Q=���Q�+���[^o1�a��n�
_잜I�s���C��|�F8�:�Ɠ�S�(A�\v/����Y�D
��� x=���<�({�ԫY�y_�F�<�2ì���Y��Y+^�]���*Fx0j�a7��c6\��CAx�*df��tS��gg�D!o�a�D�<����t�ф��P:�A��^��,���,�1KĦX�u{={q��zA:+��[G�����Uޠ���n!d���{Ei�|�����p�̙�����67k�լ�UI��^*�(kF̄x��ٳ�ZO��-�CO��G�Ll�AXUy<(e�q��b߾}f�>T"`����Xs�qF���^�Ⱥ2�%�)��N����r�7�tK:|͵��. !� C:1f}s#=������3v��"jʑh�bS��Mx>:x�]oK���1}	���3��z�����S'ғO<�^y�%{�݌&ڨ|ȋN��]����nK�v@���h1B0d�V>�*���/ٗ07�Wm�4�mF�ő��D�ګ� �%���]�w�1�c���M�\·���佚$������������?~�P�|�^o��b�;���a��/�X���*.	F���<`T̢t(��6\�@^��D_<(Ō�[Q��(~���x;��a�iϔHQxi��(My�ا+��f?�om{�Q���Fh �j���>���&)�}���A��a�%{�BgE~��B���&R<��!;��m���	x��G�e��� �!mC���GFˎY��!G�9��r������<n������={v���م���!�)]���������Q��x�ռ	Θ�V�0��L�9�22,�%�"��8hpFӖ�4Ι�l�0@�a�K\D��,a�A(�F�k3�(�f�rGt�<��o��%�6��>�9��3�ʆi�I}��C!�6`r4��hGD�Ν�6d,�d�����h��������z�`�u���no���AThuS_ԡ�l� mue����������p���"�J�ƚ4��@��4K�`CH�g�\k�ê ��2\��/)���*� ��'��'�w����=�a3'H�,�y�V��������.����Kb3�)h��ȉV(�#�6��ɛ����kۆW�%�S�Pz(�R��W$.�T�����,A؄IHl�э�@��I6�3����'>4�5�g����A��"�*:#v��<2���W><���	K�VU�J4�z]���G�Ñ�ȶ�!�t��;�Y.�t�(/�b��Ǉ�u�a��+),�d�-Ͳ�7M�1x%3 ��v�ߚy>���d b��Z�s�芤s�q��"���,��@��0t�ǌ��<|Όóa\ixSh�x��$%[Cn&G�������e��+�[�CX�,r�,/<���]��	C���9��-0S����$Rt��*����z)����v5΂��������O��1�.(�G���d�
n ,]0������R�=�.H���I1��VU�����e
�Ak&��``���0�� e�}�.�[ẻʸ�G#���g�<�̙e�A�:��m��ձ����H�I��p5ޑ0n�4��E���*p�p)H�|��`O�E��<y�B[��vH�a}��N�R̆�^�� �'�p1!�!��^~�S�ǌC��lb�T�@9�V�R���:ڠ��g^p�8h��T1��a�V�9��|Z@^~e����~�R�`>��5�y|��k ud�:�J��ˁ�O�ZȊ��s�x�8U7��֋
�,����,K\����lH�Kb0�N3��(5h��2���S{h -̣�l�a�A�X��3B�6S U7B�GP����FA�����A���a��$v�<f`L���\�� V�lg�`x0��Hfh��n�v2�����s��܏���2��U,*��.�1>��S��m�j�	jkC���O�G�<F�ق^k�9`����$Pi;��֏^}���3F>ʌ*:z�X2����=ێlڱDZ�+d�o�V�^�6����6*��62�ቂ~��K�m'�fm��,��B�@g!-����k"o7�|Q�2`G�J
�įFReG�:�� �����B0�B'���ޙ��|bFKݩ���P݀Ŕ�dk~9�K�`Ɪ���A�<�\����5�!Z���=��8\N��������o[�����h�y_)��&�L��5j����ځ��n�ϭ�MK���+�z!�a��R�:�/%�� �{�eh��<���~QC���ml޳\�����=XDS�ީ���� #����2�os�θ�H�#r	� q� `-�w���!�o\�d͍��"�0�a1`�7m���� \,�;4/������p�\.�o���Ծ2�0CY�+����<��u�O�M�U!��;R�a<aH�y#4��#��?B������MM�kfoL�NlUY�LC�`�_�ߩ��b�Q�w�0D�7-�+2��P�an������y�.�G������҅�� �V�Zy�o�7�_�����ߺ��A�Q?i��N��u�~zՌ�[&@�w^���ˁ�A[p�� ����Pv���G��8,��oD@M��e`(�'3�tr�����jA(5x�Cް���b�B�q1��q��4���6�!=_��������P�v
���7���N����=�g;:Ô�}�<��y*��B(}������Aw�y������ ���$���]	�
��P�Ɣ������0��uF��
�U�������+�X}�c��٠FF5��냘�3^)ZW���9�Ы:�5�����aDyC˟�F�8���� ����}�
�~�_�G��� ۔�t1��0�8�� �y�b]-��H���jS�Z��ԥh�\��n�uB/�;���n���y�n�6
Zy��!�B�4���F�(s)�_/lGk0m��a��5��5z8��#�������c`Wx���]�����Np9<��[�;�#�n��`ؘM�\k^�q�?n��"��j�������Z�_�&@ސ��`z�á�A%ŭ��n0�v4/��y��z|-0T)Ef�B��l�D���Ac�H䋲�j������?�m����l!c|�v�3��+2���$�&�@��ow%�/y�9�#f����C�"�h���U��\�0�BY�v��[��<�F�s`��ö��0�񭮖˭n{�����zBGH<P����P0��@�G�� ���w��7�������h��nҳ#�Y��R��8�|z��K]�zvBx��?l�|[��$��K ك-2on����h|"\*v�S�b��W@@(h;C�lG#��L�w����h\
�ϑ߁���e��c@�|���9`��� �]���-����!���)@���Tf7�c���� �l�F�A��|����u��sB��(�z��Ȑ߼�b0-��E�a��_y�/Ն���	.V>W/�O���+���jE�7T�Fq�O���R��J�c\��2y��H�ϛ���A��iq���� y=��N�ڮ��0O���G� ��1��E�h{��Z��}/��|���oѨ<��.��|:���v0�u��#?��@��5�Q>u� ��by�V����<l�������7,\�L��M6��=�����|#!��۝�eE\�ȵhh��ky!q�"=`��0<���ȟ/<�y@�< ��������H��y��q>xzkϥ :"4�	��^x�{sjj���*�|C�˸��:�;��6x��y��a�|��O�������#};����<}�ߡx0ҁ��A�.=��f |]�y9���i۝G��� q���o^y�*��w�k��u��Z��>䙺�ǹm�ʥ4#�Ŋ|'"��h8�Q6/ ��&Ho�wځ�o�� ���<���w'̗��`�|Z�/��n���B�����&uK³�q����h4��b�d�TZ�O��b������h_u�#LJ��̐�VB�*�9�u�A�F�՞z��_�����*v�E |G�����3�^���|#�{�c�|T�W>�:I�Cz����m�bY4�A�F��*|aF@���ʝ��0�aбM�Nh�;�F9�x�'��B�/U���1{Ӫ�j�P�`|���A�މ��Tt��>�����ħI�"(���C��j��ʍZ�fD�[��ym0&�^ɻ���{�M���m�!�˙�B�ccc�3�����.;߮]�D�p���|S���F4�?P7���;�8�M j)�I�Rfff��sZ eaA��$���'�� y�3==mG��#e��z8�v�>�E��	z��!_���%~s���D:m��}h�s{�l�oe�l� aL�?����z����}�F��\������Ȅk�C>��C蠿EY��s� ��N"�I>��&N
��R�k6�;�*jv:�c�b�W˥�oJ �TڋbW�&&�B��0��@���(.�e������I�6brj��O��{�(5�r�P� ���DI�S�lG�b8y儡�QB��h_����vV�(��)�����՝���r�[^*j�т���~1�0���u�·�FG�o<^xBdD>x��q�s�h��-�\'��p��	�?���I ��9�Q�a���H �v�1�[�S���X�������bnZ�t>)�8����x"��L�(��1~���imm�+�s�޽ی�O�^uC�9��єŻ�����7ub�"t0h���4^�M�0>�-�xK-�ǧOc������}����m��'�N����+���!�W�6L�|7xaa�Ҡ���n�a��<!c��rYZ����O�aX�M���e	���9b��9p�έ��u��6M�tt�/�yx�R�{�����e����B����kkccbl�XlM�ۥ�b�=�n'���H^���~5F��]��9��Q�0H^.n����^JO^YYI�����}��g
�������w��izf҄�oK��eg��A:��P�Xߣ�>j����wR�������t��)�?7�+�r�-�w��=�hR���3��2��ڦ�{��_�|��ߝ8��R8�!±�_I'N�H�3S�;�iff:ի>lNHqO=�Tz��e�c��7��8��>}:=�����0���5�\cFz�ܹt�������{��/s�u����Zz��gӱcG����ő<O<�D�H�Ї�M|�~�mo��NH���	p<~�x��7�O�?�|ڻo���{ia���x�7|jtt�e��C�e�nTI�Pػ�F���h�<���cc����_�՚����_�����O?+#�E��-�u��%��4y9&����a m~~ޮ�$z�����&�a�/����vJ=S�}�oS=�����c�=f�Jܳg�!�� �~�����������MigΜ1z1FMY����q<���_�����,Ґq�V_����g>�t��Qk����6�c�u�s�Τ�_~1=����|���瞳����_�����+�?�������,0 /O�#�.--Yyx^]]��ǎ�b��'�;�&/�Q<�1)������/ӿ���>��ϧ�~�/ZV��S�����jx�ey��Ɉ\���gB�rA��F�~Rv�A1}�H�RF�!H�����w��]��;�bC �GoDp�k��k��葤34��/~����������[C�1]��_�%�5�]��ğ����7�`H�?�h����m���r��)ş<yR|��C?�CiA�����'��:g�����|�?�n{�[����G�$厅k�+Rރ鼔�*Z�?����F����#��G�#S�x�S�OX����;�u�x��4?��d�����������\>�6D"��A�>�>����OZ[O�>���qq0^�2l�F�Tdq�ϲ��=��#ֆ�����tm9��[o��|�{~S�6L	������T�76�ݟ��O�k�Y�M� Bfya��G 2���b�YX�e����Ȼ�?�A�歪j����{���v�n��F�����^���?}���������������������C�>l���Ï�p�K�����Q�N�K/���v�W��ߞ>���7�'��r��6M�dl����n#���_Ҍ��n��F���W����6/`(�K����l��Ǿ?���[4:L��������ҿ�k�f#�G?�Q�ƴ�t�{�ɧ�o��o��}�'�����Y��}����O�|z��G���7r��r`�K{�����T���3طo��7�閿����o���^b	���O}�S�?��~���#��}���x򉩇yd����i|b2�ٻWJ�G�ߺž��RA��Wk�.�{��4�ayJ��hRp�}�j��I�\{MڽgA��wf�iM{������%�Q�)���>��o������c�J��:t�<��ӯ��&	�D���+���=�kJ�}"=��#����,�o��o�����M_���d������B���|�y�4#���1�5�?�����cR,A���41>e��_4�O�xR�D�]_��cF���?��k��C4pL41���Ld�	�_���g�̟Q���l��O�^z��oZ=^ߢ.qbC7*]P/����u)���Hem����]wݍ���O��e#�5>@���/��/����������ߚ������O<i1�]w�e=����g���reeم������4gμ*ݫa�F������S2�������˔���?`�
#"�qZ3���o�Ǜ�4�\&�幈��ў={M9ē(�Voh��d���6.��.�i�![J{���ԙ��z|�������������O?��������@#������l�v���
�	@ba�2{ՑWU� #�y�M�ذ���?��J�/����[Yd�'��O��+%�6����}�2���x�-O�㻬	Ǖ 5�,E��
�R)>�Sx�Č#@��(�9�t`$7�|�	���z���&�X��G#�'N��M�5f��*B�9��V/��w(��	^����H���B���7�P��x��>��c�U�Գ��C����/ڰϝ�'�zF�13l����y�3~�-u��KG@.x@�/�	�C����/ir�YOo������ߓ��t�=�o�ūf@,� ���Cx���#�#��hM��GL��ô��j�!�h�������ޖ!��e5l���P>���(���?�G�H����!���|�G��0����0� �C�,���I�J�>4(�"0nz4q�1@L܅�^����x 1	�cp������B�;�ӆ�7���6i��Q����t˛�dF���Fh�!E��`�����M�M+�$���m���2$�ŀ�E9�E������\#/א�K{0h�W�]���=��5gxÍOB�c2%5�^�F/�w�-4�a2z:
��"0�!�ݻ_�B�)�)G�54r/xiqń�h#h�A���R��qw��믳��G^�_��P����0�!�9=�+�..�f��*�,��Q����11@��g5��x����s?���������_�o����x?��b.�#��f����	;2��0���/9�����^�'CZ���VW�ӣ�<�^y�X:���&<������bX�2w2��N�x.���PO��"7Jn6�I�񽮰�7>@�#�Ez5�A#�i�.����0>�������6�ɛ�@�O�'k]_��WL�Љ�:H�>OB@N9���c(��P(>�<�,D`X�^(�#F_x4�$���^MJP"�ߕ�5�^����� �����t)o��ƨ+"f� s@������3�����L�$�\���8F'����0 �9���1��2�ryD)���OB,H���Ɓ@J �c��4z?�fa�`Hv�7�!`b���9�co6E>�܋����,BW}�I�F��cx(���x�xP|�0�0b�(�7�����gM�:GCJ������\WL%��h�SO>��ƃ�B�M�_^Q�H��Η^y��1������U�9G���Zq;R����%�����^�6��o�F�]���Ķt�������i+���� �(1|�� ����^Z^V���5f��Pq�?�����ȓ|D�B(L*~�G~$����׬��/���;��;f(������w�"'�Y6 A	1���eS��{�,��pO m�=]f��=tO�<n^������X��;��zxJ�CEMO��%w3P.�Ȉ%�/z��A��>�)�m(���M�@��1��a�ajz"ط_�r��N�~��gu�n�Ҟk��VuL�xF�ː�0?�P�/��l[֠��?���?���`ޙ�����6l�7��(���f���~�����ȑO}����/4⼦M�n|�������~QF���Fm"���M?�?a^���ݿ�����&8�1��\�w�,���13̡(b9z9���%���+�l `������,e��5A?��`�Fy&HĜ�N�k�@��N�Ar����̑��̌1^��9}�[����1:�`�N9��OLh���m�Cΰ�L��Gg`��7#������������~��~�:+e�2�R�Ɗ�`q`GQ��?���d|���?���]�;�e�lxÍ�3��������������4�"ʏ�؏���ɟ4��ʯ���X�����#$C�5x>&���KV������J6Lb��.���Qp�-oA}�cXq-�������.x7�Q8N^����_���^��!�k,��#m(|{}e8'oЇ蓏s�#G�0R �_����C�6�¿�F}
��|�ͬ���k����c����S��_�������$�ɐ��ҿ����)���$�Ƀ�P(��a�<i,90,S�"l����4��Pf =���.�A:Ă��xS0�H�@����SF�eqE�,eI/���Ĥ�Oy����v�y�I�(�h�I���:�O�a�y�	Ry�1����4����Δ'?G���< ��������G>��ל����������������������%�9���2��?��6��YP �D <�A�]2�c�X��pF�(J)ϑt�,��F(u3��4x��PRW
�� y�[vW@Ck���~�jhX#�׌Ѯ���5�N:$�2:2�� �N�P>)�ҐխvP$�̗�C=�yrh��
 4��v�w)�����^��ޙ�n��g?��������s���~�����?���*A�!$����@����[��V�l!4�PQ0`�T:�F>���K���:�}��qQ�	�9�.� eWD�4m��ax$�~~ٽy����/�p�&vR>ʑ���d⧣��3�	�6D=x�0f�R�<a<@�Æ
���v���Eđ��'/�8�c�EJim�6�������������Z��9���7>�����/|�����Bq��#��u�o�fSf&doƒ	H'?��@ �Ȳ e��[����P?G�P��'˛��A~P�mu�+H'O�N��v��F��o:Qg�~��7@>���| o���øO��A�4�O���M�	H�,@~�D��Su�o��Nv>t���������6=���z��i^hh��εN������l�$k\�O�IǏ���fg^=�6֫����2[�X�"����w��TJ�M�m��PV ��aE@�:��t�
���r�(��mQ���]��3�ifr����@�:Q0h��@3�'�����`�,�1��C^�i�<o�h�j�Y:��Iu����>Ys^�;q�K+�ժ��xÍO��s�n#$A FA1�P �r���}y��P,�d�t�E;��tz^�#F��? H�����߼��a��#s /(�r��ߔ�6�`mSy�]�y����LN��w�C�q�8��;�emT��gk+2��`�t���N<�b�F���[��LxÍO�����HKkyOM�=�c0����CA~�z������7GҀA�q"x0 %(A���+7�����9y-� ����>|0�r�M�;�e�؉���X<��^-e1��/���J��G��L�_��@>I�-���>7 7N�����j=�����
�2Q O��;��3���L`�\So ��?�������۞{��ˠ�iP@�G㷃0�K�p2a�j�ŃnG�"�O�a��D��p�|�2�ax�%a!�Ep�a|��'&�i3��L����Y{���z���][;G�P�y�2��Z�����Mn�<>�a?�D�\�D#����S7�x�W?���;A^P�
���+�����킼�5?;�k=���	�y��g ��*K�yC@�d�C���=��cG����.��h�(��a�܉9t�H���u�Бk�}ilb��W �ʦ��P`�9��␧ފe#f�[��7���]�7��f��M���� }
����[<���n|�AڥR��׋pCȃ��	0�K��	��K�l�!�0���G��Mn�1�1gH���Ĉ��q���(�a��	���əi���^� yyD�A ���0�uo�СSpݍ#�14ʻA@��l�����O���Yȗ�7��>��w��J�X(�c�X�%�#��L\.�4ǀ��x|s�4<�
�-2���n���t��o��G�ڈ���L4x&cNe�k>[��o�*ɷ^դDm�8�@숾�λ�ayK3������ A��4f���l~�i�1�"��ȠCޠG�%�g�o��&yx��hה^*���rclLA��7������h����^��10���j��|�7�"/���n=���7�#���E®��8� G�OA^o[��(G;_{Mz���$&&������� //ʃ�Q/�-Ϲ��ق���`��V 
.{��|�τ�'����r�W,�)W�<&�*�2�7>@CBS�*N. `�0Lt~�-���:��x�A�na��@�Qax��(�� <�0��x>�/-��Q.��1R�(E��ȋgC��� 9���NG4�b��@��ʀ�=c1r�<�`�x;��y������; ��󾿙7�Ξ�� 7@H x$@��H�EJ�$Ǣ�*[v\��);�ĥ��T�$Rd�bI)KQ���-Y�e*&�� HP$� ����{�7����wg��r3Y|�ƛ�^�>���wt�����`GH�N������f� �稻�)<T�F�7���ٰ�|��S1��oM��Jf���i� 1��P�8������:E�2�칠��7��agNl��ɓ'S�f��ȇxHK~S�E��X�b�$?�#��)g�&�8�ƥ7��y:�����O.y��YzG�HԼ3|���A#m����d:���|��Ӡ_"RG-=��q����9�*'t
<�6�������L�ɳ���#�Z�R��z#�������z�V�4�c}+e�~ld���'.Y�f_���ɣǏ�t�{~�g��$e���������O�JD���'�۱m�7��� � (P���!gw������>9���'�$�u�8����.�XǄ�C<�Y��a?	�R�ӧw}��~��_س��T*��V]r@�ؓ�����e_�I�DrNE&m߃@�@H.�b>_Ȝ>s�d.�}����M7��ի�~�ҵ��x岇�[���%K[�h��s��~�NE"�Ql������\��l�;�өc�"҉�x�v�r?����M|����'����S�ţ�^{Gk�����˗<����w�ĝM,ݻD���7}�������*:Y�[FY]�ԃlo���l"KBR��4����������ct�B� �ʆ�u�.��%���U��-_��O`�0Ȫr�d��#��I���c==����u���^���ںz����ǚŨ�
���g8+��B�'�8�n�Oݹ��ܒ�|"}~W�؀�pKKH<���twy7�x�l�UC��w��-;���,X�OO�ުt���"�?Q彭Z49��S6v�HŹa��@D
�]��HAc������֬^s��v|��v<v�M�<�K���r$Noܸ���ۿ���[���yT��!I��x�H<7�1y0�tPy�*��9�8W~��K���c̌z�PP�t:SIf|~"QsM����L��D��=�O�zܲ`u��l~ċG6�t�B� �9���7��)���w����䦛��:��E+W��\�����y���._��x"�����T-/� �-�������h2 �K��6L����;'�x�c^�,��+���|v	�yh@�'�����;�6H�!iP�\c(�11T��Q��uT��ǫW�|�+�8f���7����k_Z�`�ߝ>��k��,�`�1l�UK9�& ]�!�ہ�@Y^��t,MT�n�����H>l?$_���^���U�f|*��r��A�Od�D��m<�M�i'7�����M���6�UnW����q�'O�a��rAW��֭[7m�9Z�jU����v'��	�}HXR�UӨa�H_T?��\B�N�.�8��"��a��qɇ�uD\���ʈ�7�҅ �Q�g{��ܩ"9F;r���F�9�mFš�P���84�������%�,9�➯W�mjoo<�z��ȹ9,���ӆH<�.N�w�>G�c���_΋�;�;��cI08��(��1��g|����g0@����l杋1���}�($�I��p;�k܋E�^}�Ψ\�#��|:�o,^��ŋ�1��@K�.M�_����K�ohH��2^�U�قo����E%��*K���A9�z�D-�F�H��|�r+��i�a�%rA(�NGjR��~��%�s1�lf]8��إ�9҄�x�~J ��  F?���#���w��N��s��̾E�����E�"��`>��a�5<T~L�ɝ�4_����Og&��|r8jR�ň��{�]�z)�*m�̿Nf��'ҷ���Gl;F���IF�$d����EY�:�_�t�ϻ���MbU�իWu�w�!�aSX\ ���y̼2� �t'��G��ؼ|���3˷2R��zN��!MR~f|�'ow����u���b��k4*;L��K>�7�y$��,��Y�����:.N{������uP���|�;�E���@9��Cuhb�6���-������F P�p�J�Hq�J�$T��{;�7@�\��9�'^7f?��f�4y��u���7$R*c�`
�����~�=[����o��H�w|���j����2�����~6��=�E">�F7�-��XM�װ���x=��d0��L�[r��:t(�O���dC�Ju�#�-�cs"��_N������y:<����#�&���%U@3>��p��v��0r�:?�ʁ��@�и���M��y���}�1�K��9s�����G�+�l�H_v_�ye^����WpB ey�]���Pӣ�%�y�l�cT�nQ�}��Bn��d����w��c�-m��Χ��W��K_ל��+����G k��ٌ?<8�g��W��E*ODR7�ƶ�,d@
2��}��ӡɝ�vd���4�.t\^��E�\((�y++Ԍ�O�G|e�#kĐ<��$���,�"�S�]�A�CH��!Ma�o��e�}�̆�����Hz�A��./�2Ij$�ޓR�a����,�|c��rH���:ruzkr��*L&�Kl=����._��7�2E"�P.d����֢�$��v�z��;1L|��l���PrirD�Df78b���4�ʞ���ά�z��U%�S��k���Z%�|��* d��7np2��7ӥ�AY�?9/]3 ��&�"��ӡj�U����Zڎ��A�oz��hH֏�g��0J�5=��U����U�����*{���@��!o�?���9������/�Kgwh��X����\�p�%�
x�P��=*��f|����K�t���Շ��ߴw�ުP�K�-:z��F�o�t8̰P���x�9^M���\�x��lޒ��*[V5#�S���1�3�<��MUķfT�,C�7�c'��3�F� :@x���;�wʨ:ō=vlы/�[*q�]�Ƨ�+ ��~�W�:_�L&͆�8N�>7��=G��xg����5)?�R3�Z.z~1S��K��in��h�Ө46�J0�V�	����$s��#G6<���?x��2ݯ�_>��^x�&I����:�͛�#u� �12�G�(�۲�rR.w|�����ɟ��-�P�T�!g|�1�h$"~�٥�\���V��L6�*KϥO���N�x�{�� g���'V�.[�]{�5���;����~��%znZv���?߱o߾�o���/_�fM�z|	�!O��, tj�ݥr ��
�4ƿ �g�9���4iF�'�����nT���ϫI�|� &���s���@8[�n5ߖݼys������{�_<���坾m��G��j��_nճ�#�{@dh�ϐ�^)�lH8�1�8׸�m��;g��������=���$�l� �d9r�	��+�z�re+-�&�*�:���Y'��!ɗ:�Gͧ�6�O$��{��{�ǣ-�/\u�䛿������s�������j�A�aI��]��W(�מ>ݻs��W���`�����6��n��7�~5��9w��p��ѹ�Q-r<���,���F��Lw᧍�w��$$�_���{��gnVeb�r�;)/
���*-28�a��)��w��=Sxo:s�y����fՋ$^~dd������ܹ�G����s��om�s4I�Å��N�I�k�T]�ɤ6���kv�޽@i�a&��Ӏ�"�P��)̘�侓v�;���Mđ?_�t�/����6G�w��K��=���?)޴샊���҇?���g����ǎ_��EP7b���z4������b��#�Ke3�۶lY'u�w�(������ Q`BR��Fݛ+�`�$��C�]944|�T�6u�mG�ݱw���ٳ罯�~p��t�ѣGH�&Odڌ#�E�lM�������mr�Y	7�&����Ym��9��O�(�j����ڵ�_�ԧ>5����R.�/��*5�ǀ���������U�p��h|$�� 8�z�Q �'�\�{����\��?�]�ݠ��FF��8p`��k�5��� %�+��ͬ
y>���Dޔ�w��j����b�,17�A3>5bQ�+��U�n���,�w|��Á�N�`�s���F� ױ{�^�]@IbE>Q�xwww���-L� ��w�y��v@� UI�\�rt]^�w���7&�>Cj0YL@��ԀE�ouur/�|�Ny�H ��X|�/�y^$j�88@G<�!%�X��
���I0v<pc��Y��N��X&O L|T��uG���
9^QN�"���oNC3>5D��U�6��J����.I�	��=r��#m����I$^__�w��!��"@X�n�y�b�ƍf?p248��9�hX�G�^}�Us���&D7�t�w�-��/�D@G Ӡ"��@�L�FG<��oډ�>��(�7���3>5R��ciI���>��Q�oC����I��֯���~�X���Ƥ�y��4�g�+��H�
9_�f>`D�j��e��k��v��iv;Eʱ9R��	�N�:�0Ӥ"��
S	��Wc�S�I�y��PG��7jx֏�֒�멗�k V;���7�]�L����<C<6*}BA8�����S�x_��W��~�oϞ��`K����6o���{K�,�k�����@�:H����k�뼛o�E�[%	8��>���}�{?`��N ؁̩4x�9eSse������Ͼ}⹳!0�C���k��:���(ͬ�"H�E���`�ۤi?X	=��Cm������������I�����@!��oH�[:���4�'�,�L&���A���xƑ{�5.G����j^mdgz$!�a�9��Eڌ�$�gP�8,H8�q{�1�l (�D�qyR� -Gܣ���L�T��&�������g_D
y+/Y��p�V��E}��[����W������g?�'����+1�1��aD���`�i�����0K �\ù��:&r$�k<�3�6&�}��.�r�#q(���8�d �8wyP��	�`x����Q����g��p�<��H�|�^��ȇ{�qyrteuq\���\�o<�8����}�ߖ-�K�/:��{ї�����֎.�w�Ĵ�ToJ�`p9&����'�@�h�q��9� �����>��|���V#]*��c�Kӕ��Hhw���b|��ǰ�|��#���)��[;H����@�`�\�ρ��x�q ��� 7xoM��p����������Vz����b�>��~}���D#Z����1\��FRH��T�(�?�aG��p��������mB�R��5�(ұp��s<��6o�|9+e�-��m���tAvݵ���[$ ��;w��]w���ޕWn��n���?����1W`l�7��<2 W�O����+�rq�^���]����)��q���Cv����U�b���y$Y߰w���?����o��HD3&�Ĩ��h*�ʅi��`�c,6�s�X�g��{��8:`r�3G������6��:K	���q��>yb��q����G��|�#��>�1��������߄����c&�J>��gL9Q�؍�I9]#S^ࢌ��)9�'�r�� A���4�x�M�o���P�/�+��aF$���G�~���^~y�V��Y���0�1�
�d��"y���eC��1�K�6t��M�������a�m����͝˦�I�A���v�hHRF+A  @E�&�x6@��r9��ĝSv6�;*s�8�?�����dlǳ�j;瀎�鯽�Z#��tk�n��Oh�Ȯ#��&gj�/���)j��Z%��,Y���I&�{V-Y���>����ҌH>5t �e����,�G�� 48L����@/���J�}�#�9G<�9�� 1�j۶m�V#m�u��wv���C�	���̌�1��|,��DA��?G�%"��8�sP�ݻw{�v�2y�,�.WWG��@�D�UK�I�)��3fȦB�͙��d�����8�#'�J�e���ӡ�$/���h�F3/"�zm,n�v��o0҅�ͽD<i�[[G�j��)���F�7sw!_��{�d��x�2�K6����������I`��`L��o���:/"p'%!G��0��'��T2���/��6�OI��bF�p�^F ����:(e��`�$n��2�T�2���l������/��{�q�~����=���?����/�����e�]������la4&�c ō���J��s� �ɼ�Q�) @��H($�N�+D3�v������?��^�M�����&1���i<#��o�2���Dr!�²����K����,h��� G� �P�LiI�K�=fV�p�3�0W�p_g���{]U�D����E�p/���4�|Q���>�@�|�rC��\^������0^|�E�p�u�o�*e޻w�w􍣦ϐ>�����H�����l�Yrx�RO���2�Ijw����:"���zժ�?��/֎�ݴi3)�)���k���j�s�\�������P��Ţ�O��Y�����E\�A>t�{��G���Gf|� Ml/fv�z^ ��3�O���h�A���f��j�T�%˽��I�a����/v�\��U���G�{;޳�[�r��]ʌK._�ԫo��^|�/���Řk֮2�H9`t4y��FN� �2��P���/��<�x /�fxS"�a�����%�s�O�	6��?z!�M���[F|?��4�^I]�x0f:)@���^M�8���_��Lz\G�������)��<HC?�9�,x饗��Cjj$.K�ٵ��$v&ia��&✵�n<��<0s�ԑ<݂V� �t��z�\\�D�x�9���#Rۥ� �S��аi�#�[i�"�t�hj������������7�q������Q?��#�K8L�wH����_��x�L�Ӏ�=�a.�w��9���4ŎT��=� x�ģ1 $�4�rp�������2d�3@�@�̼l�h̎'�)5�� �/���Vb^N �dp����q�N�3.P~����ϩ��1\w �|�@)�s�(�-��@�>>AN�P����BI������k�O~�=7���E�V��.�f|�g��k_��~1h�3p9��|N�Ø�(_�UH�$8�(�(4|Z��>g%&�b�Q�LZ��W�7	�HK�M�1�G#ɢF�!y���3X���/k��җg���q��uܕ����s�I`���L&g����$\'_��9���H\lL�uC>G�al?�K�:rN����L��pR��US��Z����[��ۻy�v	��NǢ�omݹ�3�N��$3�����������k��a�gz<�c1A4bߣD�Aa>�/����j�Tb���(G V��3��F�>`p h���i���aJ�5 �9d�x* A\��TP.�0��ە�P�Y1s�t�iऐ.����`ԓ#�9P!�LG
۵���Y)�s}���S�ԟ��>��sR�J=G�: �x�o�-7y6\~F���7��W����y�i����O~r��������� �0Ʃ]���8�nAh�j#��T�R�w�u�i<1�� �h��}<Ѱ6o�`���gL^���9��H�#�C"���� � }���cR ���x���VUy %�������Q&$`�v�&��>|ZiG����+W.7�S�|�;�3y3I�\��Lo�v}9y�G��$��%��6m���P����7}j������ߧ?��_��W�VRc^&�@�ƒ�s�*'�bh��y,�~����s�=:�L�a�
	FgRi#�h>����ۅ��ʃ9c�ej��N�X�dng��&��u���O�6��%M�fKc�$��<�h�x]B�R'P��c0@����"Y�<uu�o� (�N������:��:q8g��t٨ ~08�
F�S�o|��D�,A�:"Y�{)>ce҃o��*���c��������m��F��L�X����o��^z����0�}���ݻw�OL���9��Lo��H����x@�M���w�af>������w�kl!��QS�}�Hc J���O��h�@�QM��H�t�2��@@�ٳ�ip@u�̩��`g�k7l;��1� �g�5�8�l�;sz�1��$�RJ�:��S_R��	j�Ay>���&~.��o�$S�+�h��˽�a׮_�.���|��	+4��h�����ѳ������iSS���%����ȯ.^���/��i�糺eHLf� #ڨ��h&P�q�<�Q�	�C�nϋ{�W^�o�d@v��� N�QC4n)��(�3$u����@�.�nNq)+�?�/U: ;qhԄ��!5��*}T=�*�4��I����� Pc20|R���J
∐w������Q/-)�\l�{�P�u�z���S*�M�T.�� `�.�g\��8P���h�Ư��e��<�H$V��s3>G�qgeL3 �\���Ro�ˠ�M�a�����:�;#��/��dRc�H�Ӑ�����#��%i����琒 �����~�3�{Cz>�T�HI����݋���^B*�1=����!�8pG<G�N��)��R~:uÁ���3B�Q�Jl���%~:���Ư����⍬�����ͨ�#�� �	h*����6�SZ����xS��	�=�ޱ7O��ׇ���ߨ�@���`U;:*���%�hP@���"��d��*�$���%�L��>�������t <�z)Df.dJ����5lx� �lfl�c�/�EA�yhB��3I�Gd��������s��;y�W6�a��}�I�W5;��P>�M,w,���}_""�k�5(� ��B�z�_99Ra���O�v�����`<B�?�z��R����~��	d�f�9iC~�1~�&ĨT�<א�HI$,R�gS�� M����ᣦ<Hi�Əg 6�K��r�h�����~�<); �/8K�������6��}u���8���;]�fXu�=�1Ud��T� �ܹfT `3A�H�!p�M&�C4$�h���C���� 9�"�Ni�@F������5�7�G6��4��β�ä��� ء�w� (��.ã��9��Z$��Јʉ1��l�9��3�@����Tj�+o^�<��9ՇN������9���'��<O!�_�RU�"�WN���?u@qՠ�S���Y��) ��;�����k0 F*��J��?��X����ˣR��!J���q �q���G���H��wHزKbP'�	~s?�N�
���	)H>t���6vZ�H�4m��	��$M݈�}ҍJݓ׌箴��Ĥ�	ұGs0䮝�Jqt��'�f|b�Ķ��
�h��T�8�c4q $���~w��pL��1�&��^dՉCx���˦3����iD�9u�ţÒp1c��Q2�G�H��GBK��J/"�2f.�
�N��=���uI/��h���� jg:b���^2e5)l�Hz<��<���x�د�b���_T���^��6mG<�Ε_H�UH�v��1��9��T����E �|� *�I/BL`b��eO��Cz����4 �U�w�Α�ߦF�K^.p�ܨ�sf��6��%	iq�r8g�8�@BY �/6X:Ec��0��S}x� �K�Q?���/_�9�n�N�Ʒd܉gTm�Z�JB�3�S6.rDJs4�T�Ai;�v&]�ccD]M����@��r[ѵ��_�] !�0��*ȑs� 8w�9�w�c��%.y��6d�eb���(�` �a�Q�n�C6+ȃs��4��u�!Xu�����(}Җ5j�F�SePa vHR�t)�]Ulm1lM�	f\�l�z��ժ��Fz!��[|v�@١�_�Б�]C�\}X�C�&�u2�W�	�OӡEa������N��k3>1���b5_"��0��h,��5���8��#��1a<��\�����Xy�g̫����R/)�*O�I2CF�߇�|��S����s
�ϑ>�<�Z[����^w�<o^G�7n����c� �[X�b�#Rv�*σ�1�h���ލ[��n�z��庫����}�F���eRXv��y������Xl��"W���=3N\�h���#*�*�AE!��@Cܹ���d��xFsD�p��'J��b!�-_���r��j�����[�2}� ��4:�|D���d�!�vA��Xҥ�����+���~����[��w����9-�i�-5 cm!k'L'��G�ކ�H�(>�綷z�ٱ����1�w>~���Ȼ��[��4m���qN�)��Q�*)D�������%s�����u8�c�>�L�D\'0��ŧF�ۤ��
�8*M�H8'8�PyFr�"M��sNZ�a�o�2��X׭_����z��6���ۻ����Rw�
� ([�ĒG�e Y*i�<p\�sJ��uk����^������#޲�f�{�|����	��l	���X�+ݒ$FZ�c���՛7I�]�m����k��.Z`�&�0�=Oz�g��R���:8"�t���� ?9w��?C܋�c�X<�hK0�p�Qɧ�����x�w$� �]�i7��2&^�t˕r�N����6�-Z��m��ro��W�W�_��8"4j���9�g9�(�P�������-�VY�.�����yޜ�fy��n%�gȇNa�����O�+q���H]!�$���6�x��:��>�5�u�fkʪz�e5޷@X�Qn���0qʃ#W���n�d�F,���k|*56���B�`�pQq~�7�c�#���h�����$��A��~�J�Ʉ����%��jH�B�J~�]��*ϳ�,�͋AH������;=j'�l���Ƃ
ba*����"+O�ZP�����K�>�*/���Ǜ'�{o>�z��L�I�K�������(�y�c�H�o��2uE�s�����T6�6�)*���0*�L�P�X����i���2�0�
�f` �Ό��4���:$s�h%#�J&�^ϛǽ�o�F������q�Ō�7�<�y섗�X�S����I0p$_*Y|7���U���|V`R��L����;��=�:�ɇ4LGS��3�e}�eeP������{��� 8N <�nO�w��1����^��^/��zu<'�3$��&"�u-�N��$������p����1UUP}�c��\�OP�Km���Ţ�q6�K���L3>K�*�2ڪQkSX����ʥ����G빘l��� ��\�0��T���� �����>3�q��p*�:�C.SSvٮ�@C�v�L���-m���P9�3Fݹ�Z{��0L����P'��	�N�Ho:'�żt�sx�H��9��e�E8V���$	��Qc��u���	�*��_������s&����S�Y�Cc0u
�[�c���J���M�Q��)j�:Bg�E�q0�^��$�܅d]�̆���.3o�1�Ac�H�>�R���7Җt�v�=T�[.( j����Z@���8��ⱄ�
l�2s�Cހ~��%}�_�H{,=�� �=
��-yn�ǳ��PnV�p.��ۖ�@�)���P9$ʅ7�#t"��r�L��ۂ��Uy3�Ʊ�"�sۇ�XU�ÂX,�min9���t@Y|_��T"�2���(���v�I��0�߆��ƀ,-@`���`���0��}T�5�գ%��X ܈z��0�Xi2j�u��~*-t�$��,� ��=ǵ\I�y����\V��;&3�����bj���z�lu0I�(6�BL�0�N�^3��7��ܠ�1:V���t5ľ�ʯ�_����z���7׀!y�eu8�rD��x�K��(�,->�S�tF�$Wft4���A?���������4,>�$�#��������6��А8��R�\�niiy�����_/�olZvp�UY.� }�߼�_���8x��Uj|�0�Ӱ�����C��q������l�������$�Mި�&Lu!u�l��ݰu�idԖ��R}��{��}^J�ၺ�[��(�r��7�#�El�ʜ���^ /w�3�K��+�m�7O�x}����/P?�;�MhHr*gJN8�g���0~���
�!b����]ު���R�4���%���/������*�:Hj�ҥ=��������é�t 3����z4�GU�|*����;5W �m*�)�^�p�˗/y���+-��p!�΄�L���f���D���-��ߗ���U�7s� �Q�����4��:�㚓<�VǴRG��+7�~�?��n1���}�o�~�;�ެ^�%�f��<*lѢn��+7z�O�5�2u�#j�С#�(����L6xi�EY��kt�ҥovtt��3�t���k�?~`P��$��e�d����a̰! ��sRÃf]��D^?r�M-g���~}��������W^���G�r���M��u�/H[o��No��ETE�C�.�ۀ��=\.L��\  ��t�˷�r˷��ǲ��  4IDAT::Z���pNX+ȶ�%�1�������N��X�����MM�Yߟ��7oj�4� /�p��%p�v0&ӌ������+_��_��R��D%�!5(��h�Mh�y�OjBNSl�Ӛ�䒕����KW_}�+�h�����~�����;�T�CG�:�u��f� �S����V�CJ>�'�'	��ЪU��}������������g���?��'?j����mj0�;����ө�Ț5��Ɔd�i<�hԻ��2N���V.^����}���˗?��{���M7^��ҥ�v�>����~����?~������X</��/ė�X�_0oA� ?�o�H������~���A�،@�R]����7n���~�_n�z��*{�h�����|��駟�T�omkk+��m���6E� �IL�̞�ȗ�Xb_����{6o����_ޣ�?��3˾����|�?����n�̰�e~���UWmD�$� ^�Db)y�#INyg[Zچ�<��\������=߾��Y�vɛ���Z�СC�d2���ݻ�D����IU"~�U�s��@��-�����g������I�c�3s�d�ɫ7_�Ķ�m{�ŗ�m��ȮG�����{y��R�M1%#U���ȄXs�رUr:�dn��u��\w�Cr O$��B~h��>9:wN���u������i�Q�nҌ�z�Gd�F�?���s�?*:����$LQR�(��mۆ� ��ynz��'�?�Ѓ�O��
���2���A6�7ԝ�9~�����#����ڿd�ҧ�GF��������áP���ի�V�Xq��K/3�?��Ot�۷�-�)�7�4�3##�$���?sӳ�<��`./y��^w��ol�p�S͉���SZj=hi�O�_�e@���l���jo�����_�M>�̳�=�ē�F��J�S-���{>}��۟յ3���j�f|�4��D��ii��Mx�Tt(��:���z����Rkr�#�6o���;��Ayu��d����ʕ+/h������_���������̙�k�-2�����{��G?z���g�	�/���k��'?�l_o�FlaI����������ֽ������P�;M���������W�x�;v������tX�ď��h|�yN����GV���g���
<H�P<�e]a,���p($�+���P2�"�X,I$�~4���G���Gj����TI&�|.�
q5\4��d��s|��<s�Q�i�HT	g�����$�3����2��a��]��w"ǧej�f�򣣑\�OȖg�;,�@�$	�Ҏ<Ϗ�紴��~�mm��`�E݊)D9%��WD��X]���MeO�'�E�W+����'���=�[-�Q��ʥ�ҷ���
��*R�%ba��T\;�:�l�jcn3A�|�C�����p$�0�R��M��@��)�S_��I�%(!y�ъ�����
�S��<�<�z��3M�|~]]�H��L����
~��y�ڳ�=.�I��!�Ǵ�Q�n�(�NWeD�P3�x(i#�y�`�l�:����B>�c0�P$���[���F#�@bTG�N�C��?<<\�,��f���(��^1�My,i�]�}��
����f�z,ʃ,�yT[)ʴI�c5#k�$`��Q��F�i��	o��*.�LѬ_.�-�����	���E`��Y3+�*���=+%u���`KR�R�kxЬ��jN��5$� ���'` �0%�z�eXՙ�R9�,,�2�OeG���I�w�f�Fd����0�3xe��T܈����a.��҉��0X2��3��]zFm�Z�b��:-`�ӈ fDD�*� R�E��G�$3'U�ROi����Ǻ�i:�P�gGMV�J2�2�yǫJ�90���Պ	 �nm���M��Y>�����ʤ�x��P��+�w2�������`��MsD�Ir3�X�SkЬ_D�!_�V0a
�������*��))0�B,V��30���㬃(�kD
�(/�W�m8���E_�p�O�g����/902��o�a;���F�C8�x^��C�&��_T��D�Fͫ�%�ɗ����s�t��2�ER� �VE�a�I�R�����ڕ�6�:��D�`���|���%#ib�G�A��G��H>l=QN��M=J�j�f%��i����8gΜ�@8�bŊ�AD"Ey�|��|c�(�nWDr��!M�Q���n�Y�v�*�A�2g���UQ��p8�+��J7�P��G�$�T^^�6ӂ�}`ͮb�f�X�f�Xd��~
������p��+�v}y��x�Af3&p ��HJ9)͂�>����ە5�~g��c]/`)�y�zpp(�JשQ+nD��bT ����A�ޭ�tb����B�s��r|�DH>6�@�!=dě�jx� �mg�� �-(��tU�e��l��>�)��c5ۆ�P�Y�$�aW�l�o�(��6cx%�p ��lw����e_!�H�(��G�2���_ �
��f/�'��E�"�bvE�b��bQ�*f2�T:�p�U�
8X>%�gU��#�֨|.��Z!k#ü��p���Z���Bg�6��I�_��%�U!:M�'��[��E�WS
���D|�	�bq���X�y^��ds��*�v�kDcՙ�P�,����>��jzv�u�S�	x��NR��#��|��>��A�t
�peJq�����KI�wO���Z�]�4��W(,E2���b�6��`�-V }�e���l�*�#�t�K�B\"C��"�:��ZL�<�� �cg� v�p�Ng2�B!�f>U�@�N����0P^�]s4����Po��@��v���M;�hC��͢O�����l��|��g9H|V�� 6�k5;�6��'iQ��Ǭ��#���B(j�0�|�c�	͛��d]��P��b������}c�:��t��/z��Bj�b���S�k�{~�:+Ob�@�4ľ�|��3u��Ƙ>mڴ��݌�'���Sq�f�pց/����##���A�i�3��S`K���� ����I�V5�2$_N���0��:{�]�|�B|~6�Q0/��C^("�:�ܥ@��AN���g2	��|�D�FQ�|ؔ �1�R���Y>��H����2�V����iR8, ��/�o7_�9��U>+M�3�<������vk�b�|"e��&�x�B�W'U,A��p�ɵX�~��7��ď=Z>#�t�b�
tH?�����\�(%�lxp(4:<�g�qɕ���D�� �#�EVE5*pg����fqD�Ҭ_2\Whok���(�mo���)&�+����y��`��1Y��t��7-)��"���GbźX�J"f�f�F��b�A�|!T,� Wː�x'+_,��)5��[__�f��S�W'{5O�?���T&-�.�ݚ�|����K�1(�s̛��+&��E�~����P�j�)&�#&����dҩh&��8�RK�t`n����y��*�$�%��'ЙY� �Y)Be$�Ti�ޮl�T(��F2A��%�Oj�*���8�My^w�v�A<+�6[f?� �K�U�s�a9�)'kxC8d�I�&�:��0V�e�/�����6��)��s���9H�R�.VK�F0��a����H���oVJ>U�� ���1>Y^�L�il�E���}���)�D�J��c�^"��x�3A�|f�����oo�҈AP(�$�p:��H��3�W�]�- m$����y�m���ڣY���Ʉ�!u	��:���{���/��x�FKw+���h8W����!|o��Y>$�j-�1F�Ћ�HU�+�p��Q^i4+��ɤ���KQ*�8�O}�Y�tZ>���Eo�� &uv1i4ZZ�\�eO��3�#s��1ۯ���@IU�O���G�h�7؊�E�cs|�B�|>���� �UjLV�ŤK'�N�$M0����|���9�"�b{���X>����yE�� s��l2fFrx��P��k��(��L1�ͦ>���J�Ϋ�真��0���G�S�h<���n��:���X� �/��p�|�PV�z������R��H4*��� Te���)9:o^��u�ޠ�?#ۯjj�ݦY�px4KĎ455omm}����P,)ݮ�d�v/�����w-X����8)m^�����yj��m�z�οܱ�=_�|�U��>�L�v�Qͺ�ӥ]�vE_y��ա �*QW�(?w�^ٸe��R�����_�����{zN�:uꔌ����H�V�#l���}������ŭ[O��>d����:�A ����Q�̋��s�^:\�U�M�����E��esΌ�BWVx�"]�����/�Zձ����    IEND�B`�PK   �r�X�&�}[  y`  /   images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.png��W���x��,@���$$��[pw'h� xpww����]w���{��p�sf�L�tWwu�S�]���(�P@ ����2s��{����[�<�[��)Z���@tq&����醌����Q�ܕ�ã����0��Ќ�P"��b``�E��X����t��a9�檗�����EV�����*f7M�?!��ģ��JHH�`�s��m+�>=,?��8�B�ybѣo�h�I����7�.5.��}7�O�3�����1�]��fPz���	l5\B�zB���Ǡ�9�WQ���t��ԇ�t�D���=$9���y?����K=�`�?y.��d�bh�h�� ��;|4��e44Z7���A!Ɂ��Lс3N���R����BS����d�����_^��Fe�v�����t<����)^�"��y��(�N�Eİ �7�R���h@��`�(
��@�� Ё!ğ8��(	/�e$�A�]wb���?d)-g���#���(Dr�����C�G���!I�_��������{'{sK��.�f���P��z�>�7�Pz/x}�^�ʧ����f+%O)%�.V�>�9y 8�o�Y�ڢ�d4q}�o����V��؂g`�`࿘��u����_*�/M�ܛ�C�M��T��0=��������,�.^��_�������8&3E���1]����ߤaV*宣�K�W����?��P��|����������gi�j��fJeSk�$uQ��h�/ڳǠ��S���+M�x��}BM�9�+��rE�4dMӌ�����b�hp@���/fg�����Njy�|W"D��=P� �LC��˟@2b��+�U��=L;S[�1}?�	�c�'�z�ײn��Q��I�g���)�GD�!����3KWEc��Ǝ�YXG����w�W���qO�t���?�z,�����=#�Mp�����9Iq�����]fn�����\QQ8қU��X-�?�瞭���ܷ�Y�}x0���]���Y�c�����MY�W��Q����G�E\ж�aL��f�y(�3�_������ţ����6����)A�X�֕z�ΉJ+a��©�����\l���f:-��¹�/t ���'"�vy5��S��Y��u�èh�z��x�ۣ�ni{0xq�ʇ�|��_#[���%����*��5� ѬXX�'����K0y &�>�NTm��Q�׋E��j�@�	�����z�f7�*�������i�ǐ��	z�M��)+.���"}Ƙ�s��̥�b���93�R�R /�y5R��w�>�v������Fdt���v8���ډJ$J�ݜ��t�+�~�?<��la��綖Kц���x��+��0Z;H�fp�;����7.�c�sϋ����?L4j�ctҲՊB�뚚�&�n~��/H�X�A�uM�Y�����5�W���a奫�r��E��泑�'�'CR���:N^��#7�2�d&�o�ȩʓ��_���ne������;]V�	�%�R=r�G%N�UH	�|:��}�$�$SX9\:�H\�.)ah*-Ywkݸ��l7��TrCnElN9�����
��xwy�����=����$�a�V2?�I���)��5V��'<<'EI�I���%���-cO3:�u*b҈�Kl9�@V[�~%M���0`r�b$a�k�G�V����;-����m�'�{����6H��ca)��rw�p]�s'%���R�զ�ţ�L�L��Iծ���_�me$-:���y�'N|�ޔ /�B����(������\���y�I�f�f�~�ٸ�(ka��o�e�����{�)T�,K}!Q��`@6p���5A�`�҇��P_�3/A��8yZ,,,.1FF�Б}��'?�-_arFF��#��k\����~y�STf(JKI��efe�zQ<o��F8���>�!�lU�{�)�p�w���,.vj|?�!܉)_�1���ϼ��+{HQ�W�gmq��@WB�`aVN�)A,��<�:�^�Y��CJ,޸��o(ǜ ů��gwm�@���8Xt:U�.�3/_V�X@Bs���8�&�3�`^?�k�of�Z�0���%��2IL�P�������d�*�5�-M=���m�D��I@�)4�
�wQv".#(t"���k���R��,�WR�	 �ϓGEe%P=|��^;��_I+[kRk����J~��(�:I ����|8��d��%���z2=1�+�u���k!�p�P/>�/#�e�4�������5��D��t��*ɟ���8L�WD0�OD�(ɀ�6�a]V*�,_�r�קbC4�\ $�1�xJ,SR�r��z���oTgdS�[���C���m�:-���5�t��I
�KͿBʜ^%�*��'�����4f���Q(`���u
hR\.
���쳜��dMV�#�������IW=��x��1�ʐ�ߢ��3�����B�%L�D��!4�0+M��f�3���o��&x��-����Tl��d2��%E��`W걆���	�ε�O}�!9b��7���ʷ5���$˛j.�����K�8�j����#�psJ�{"��<|��[�v̆[�mIR+�?v��psL"��kDs�X��ݕ���)����2�_0E���c�3��Ȫ���ϧ����t;�	
�UUUlbb���n�F
66,�jA���IL]N���ē�E���((s�ak,)d o�~��oR��}�Ku=<��1��Y��t����K;y�V"(���n>��0��W+���,�P���sB.+ܚv�iND7J�M����w�r3����'{
���k�����-���4�j�cm\|\Ѿ�o�s(��+�cz;�7�������ⶳGԡ�5̙�~����@8�.c��m�� XE]m��� �0��a>�7}eY�՛ł'�äa�.<�L��ۄNm}.���0s������O�TUL��#�\�������.'z�	�:ڽa����H���x:N���w�ng�4���$�S����',x@���2m�]ەt�QO�ϧ��zkZ������ HS�f���`�eg_�;��l&F�� ��۪�� 0�A~�����{8ܙ%I�[��������灚��|��<��':�N��o��P�4L�Q�z�������4�c.�{6�?�2 ��U�Tv_�&y��v�G	?����W���4�apP;A��U�4�K$�ԧBG7�%[��r�6k�n4l4��i����=���d�0�����V���`���C��s)I�=�%/�4�u�9H���Q����'�,W��ЮY�B^ī܀��;��@��T烌(�7���v���98��Zݾ��1�����78HEC�xR�����J��	E'��=����Ϫ@*�^/+�:*��-�C������r�(�*�~3鄖>{�q�/���f�H�ܐyV]/�����ްd7��r�ߦ��0 �jfjn<:_���2CYV��Ç]V�v��+t��%s��k
/�w�{&[�s\4�)A�k�=�v���-7�#7DW�������"��yZ �2n����Ir_�ʗC��62B�̘�<�t~_�����Q�l$Ȏ����%>�=v��TpZDD���M�Y-�IF�/�pq�{Y���<���s�OW��Ef��iΉN���ߥH�:�0���(�8�n�5;�����;w�+�O�e:OG����\{�B��S��h8B�ޅK��NC?:=\K�{�����x�?#U9l|^}��r��'��c��)�=�Y��F"�쩅��h�n�x�ﱿ���ܼ��B��˧�pPx�����C�!��Gx��|�%���5Uq���pH��}*��^�{V��cq៞=����U>9��e�~�	��b�u2�++��pR�ȼ�굺�9J�ޞZdn��w��g�C����R�sB�x)�vb��/WS�֘Em?`�r,���]�<��C��H%�>�b��)�13tɰt�?}�2���x��iz��V;R}�s���7���&g?)�]�>^�>����c�����X6������I~�I�%���5EA�N���l�b���ͪ�\�N+>kr� 77���H=!��<���,�-0ߕ��D��II���"aK[|�|�3�e�_��z�;�hO���a[~���`�Lb��e6#H����M�M���*Hd��.^�$`�8�{=�r�w��K�~�y�b�x��>o\>l�{m�`/�y-w)�z)�ym����8I��N����[ �:x/�=<Ui~��.��*gM�E�77��El?x��{�&&nظ`X�iؠi��n_ن�8�p���n�t�Ab��K�Pd\;����.��o���BU� Y�%F��Bp&>�ß���]����k�k����ֵ�}�APy����5���K�M�K��k���r��jIy(C��EO��N�/��+��sU���ؔ�¸������Z�x�<A��u����d��:����t�`����zC�W��_e�.���������vY�S23cA�r����(hi�ظu��뒦/�T�չ�Z�M?ub�F�(n�f�-�u��>��f'L�������0��:����d����!�J"F����g��ɜǒ��9�*�a�2�F���������d||��>��hd����T��cw��J?~\�ή�Y��no�j2���dd`�n�>R~mH��D�ݦo�>?0�#�����c��E�jR��� X��<xkpE�fd��
��b=*�2 a�SW'@#��E�������|m��R~L.D��8��\��ݿ�Zj����'����ic�����'�B�5�% ����0���[�΅ʒ��Җ�3�I�R�R�_����)8��LLK�\����o�!�����~���x���C���?	E#z~��*�f�.ɫÕO*�q��ɡ�]4�+)j�n	�ܪ;/������g1e�I��Ӣ	@����n���v���}f!S��G,��"�\V�[��X�|
fa��"�L#K(i�X���|��S���r���^������G��R(���O���moMR��t�Z�8n>����U�!¯﹣�v7��76I���x�y_�B�������n���>?��|	J�+č��YSF!��8�|(��|f�C�V��d>�{�U�w(�xx�
�ď*�i��=Ճ���,��1B7�}|$������8%�A�G���j?�KȥBIy^���m�7�-.�(���EA3��3Ӭ��ot���m���Ә�N'&�2��ڣ�e~ge�'oY��/%���$t��j:�Y3ꉠ}�F��殺!��`��xg����ua6���T���w��j�2��KX�Rh8��2Yn�F�Ie8y��2_�&/))�R]�N,��M� *�� ���v{68?i=5�nD�2��ed�:�'3�h#"ƻpz�Bと}�R!&�����'4��[�oڮMJ�����������b��$?�_X�78���؋�U�D*�H$ǁ���I_�Dz�ɳ������]\\�L�z�����̒,eL�s���ꏈ�^K�G�L�?��.��a����贼�6��z�"��\�ęq^�_�*��q�h��{�c{����y�
q/mw���0��2w*�`��Ĕ�/ Q�4�����;M[
��L!X���kt��k��
�,	������D�qh�?4���r1�U<��֘썫�M��d�q`�+o�����4�3'^��S��$�vUGGG&9���Ե�`����_B`�����
�V��@C=��d@A�mk=�:i�ޙ���A%�oe���^�c��~_T}q$�B���".�g�de{��qX���.�􎏅{(~�<����r��ŢǴ�?L	��7��C�fo/,c��R���&kπw�o�ӿM[P߾Ϥ/���宥34N#�Me�O����l���O�MFe��z�Aڊ�G���p\H$��g ��4��[&�D���5)=�gRS3��}�
�f�fn�V�����T������bꞘX�.�g���^�����$2G;���M���
��`JJj3����2{QeU?�rS���fL�Z\�����tfV5��	�wk
"s�I��Ѳ#n2�_S&c;?0��{�6�}(��r�KZ���H�|;��& �����kdw�6��>�tC��-Kwк��R��˵���v�VzWhi�џ$^҉�	�:��l�s��am�ߞ��Cn4�	!�J]�����X�'Zī_��>�a�����zQª¸9�����B/n�Y^��.>��������4��� JBq���P9�W��+���'$�J�Z�T�L=�J�2B��B�x[7��_��/v�aTv~�K|闦k�g2��W���Z���صh�T�{m���:ָ=�/��W�%x�dP#G�d��(��4�K[�%���}�W�Tg.��� ��|<m�����P����"�y�9BIy1�s�g�Hv�v];,��n[���D��7X���?vi3��b��A����>_��9�ȸP�#�:8ty������/�+:�g^�~e'k�ħ"v���Z�����Z��{j�#���_���
�d�wJ�Q���N;�F*��*`S�"&��V����{�y��V�Hs�y�b�8\��~/7V���o*�֎j6v#g�{�#,�E�,��-��d�K7
�8nFA(�k�]%��TA������	����E�ʭ���Z��ʦi�D}/df��vB0RǮa�qw.�rx�pZݹbp`��<�Xx���I@�"W���b0;}�n��ZA䅤q���fM���~"onb�p�K���a��#����V�Ksj��l�Y�W�cBw���!ʋ6�\���3[��������|�}�ƃ[+)zP��,�UC�R�?9ϲ��=�g9�Rμ�|���@B>'ܚ�������EM��У���*���Gk��-�U��7��MwiF�K�����*,��ka` p\��;ط#n3�^�̗����D3/�%'�e����&�*�&�v=TWm��`���<_f�����֣L���fH*]u�%���tj��ҨԗRP����e&p;��p=A+V�2z�&��56���cf&xI��C�%?c�A�<N3�7�ԸEHij�R +��@s�)(`����,q.lؚ�E�*�۠��[����A@�����s;Rh ����d�x�g-mup��o��h�N8󜳿e-��~�pvlv�JL��aI�~��+aӿ(	3O�I�!3�,Q����#Qp1�;VW;4��}�(��O�Ϭ�z�/�,/O�|�i��%,���h��ƐF��>N��@8�C� �@+* #�\ ��sz�%����Ca?�����]���Ȫl�0�
M6�P��uϐRn�e�A'�W��B����څ�U� >�,䝚ʕ�=�	P�yO(h:?�]�\�@��zb����Se@Iy�y��yh%��SR���_:I=�(kl�Q���\8Ԅ~^�g씈�Q�v��_����AeL ���i|��d�c��ijfƣ"��/b���j�������(���{��q���Vl����FiG�&!��{��s���en�Տ)T���hZ;f�Z���ӵ�w��
	3�"*��l���22��)̫S�gѣi\s,��vAM��U#�r+r�,cT[e5�5��"��&����js)��ǓQk�Ro���h�6�>d�{d��T9�b�˒uڔ�1[���Qr��y�t|��e�3�5��l.����kA�޷{A�}W��}m7��}�;_�î�1PcE��.�k\0��Z�	+'h[�'��"w��O�^��3�#b&�t֗�Ǆ;&�*�H��'�]���i������K�C����umm'M �\�M�3.�%�G��2XΑ������H虙�d;`�[�Gq+�п'B�fk�p ,[�u��~PU�ɩ�ڍTc���eq�ys��9=n@����`�S� ��-ڎ͞�s|��9�)o�` 3X������ܺnG���;��RJ���ݧ��8���[;���+t�[�SR��)�������%w���ݜ,�=��@�����3�j���-�x��6�.8��4ᤎ%,�4f�=��30[�	�g*<?�����ɱ���UDw�Ɔ龠f��Rѹ!�Pg&�hg�����xFg���V75"�Y>�->���Ѧ\�ݑp�\�������Et�R�h"���:���3E�͑�ne��c�g���4�Au���˼,��-zc��429��/1"FA>���JX�����iX�n�]��g�����E�I�w����#"�?�yYY���t�H��u�K���sz@J����=�{Mm%~���lg��I��5݆�%Ɗ�0�3��FcI��1�`Y����Z����2��b��y'~;G�4I��[��eU������׎Z�G�*V\e�zM�s����^�!T�Y?��c����_q_���Z�) ��村���!?���w<���S��t��G�9�rc0s�$�5a�彐��|̯���?�vC������m�<��6v(��ZҐ�:��~K�����>�i�+�Ҿ"E!�$��Q��A���r�|����Ö��:��7��K�����Ճ�P�eWa?׽�u���Sޜ���bL����I�ZUL�y����\��e�۹�"�p��`���x�l�'�K�}!���Na�� x��Sn׋j����BQa�y��V��1_tbn;�A�l��z�����T�zM��0����¾^�2��B/M�8��7��f���n�h�m�tC��c:�L�.��͒��5�',���/w��}���%́�����MO�Kl&�œڬ� ���s���K��\Ee� �������+�k�RU1�A}y��~��M�O��:.h֡^l�!�����[���s}��/�Znv�vWܐ>�Z&{��.����)m�!���_��:�S+j���>���f*ii-<V�(Z�L>n$u�h`��5�A�GD1s�����z5�o��!C�����n��7'+�D0�\č�~�����$"tkpE���:�l��#e�w�p�is?��i(��a�?��8�%$З�%n���"�ܔ��Š�\Re&��Bj2�?���['2�\z��o_������P��t�}���#0�m����J}�"�_���c*ӦF���s�t�ڎ�=�.Ǳq1��KM`��j'��9�"��]E�J�迬��a���3[�ˆ���%�U8��|.B�
j�F폼�e��zk�(;����쪢"=e��BK�F�k)�������_	\c���B3�/·�bM�x��5mo{�_�b��KK�$��\�zHaT��& �P���9����Y�@�kZEE�	CT]?����u� �c"����������I�#`�U�Gd�R:םqm�z*�(��H��QaM�ڮ��2�r� �I>��;\����aGo��cf�d������l��t�k����!m�]3@���mM?U�DH��BF� 	7�wqOD���@�:�w1?��g<��;��%�㚰/�)D�*�#RI_�Fq�?lQN��T���,F�p%A�.l�
�~^á��j���gɵ_�q>���b�%8؝���@,*�H�
W���]]b�����3���Z�	=EK�"��9xk����ۖ�����r?�AYI	K]�3�g5W�F��Z�ZZ��gypE#��(!��=}(���gX~��&�/_�.)�N;ol�ޖ�رk9<��Q��4���N�	��Z���t>5��|�m�W�b!�`.g=3V
���3�z�c�_۽͈K�Zbw��2h�u�4�P��,�V�m��h����t�+]Б�K���� ��T3�|�_��������ݞ�> �$��3qm��-�p�~ 0���E8m%&/�C/4�uM�g��5ب7��=�ưZ�g\�Q��iV�٢E�im1
��NN_�}{��!��t�gy��j[5����v�E�X�ڲ���#��LH�*�zw�Iҕ����������$\�h�5Pn֔����%�E�ʢ~q��k�>ߒӠr/�	Cq�x�m�俙t�q>��M.�r���eu��LS�v/A\>j������2X&�����,{0dOy�#�oY��UJJ��-���q�{�F��CۤE�|YB�o����:�g8����������!�Y�>���c޺����_p0�0�B�0�� �H_.q�-��NP�qɾ��c�-��wD
6���.e����m�R"9aa�0�����IP�ԗB�|`�1��(��ZD�v�ߚ*�Z\>u�=ah�kq?]��'��=��&��Ňg�@�>Zح�JEl�,��@KK�*��h2�s�����eU��~�o{��e��ȭ������T��w�����qTjR#�7�$P	�b��{�dLwU��IS�ݵ:K�4{�D�l��?U�K��l���g��A1�a�D�RK�N�369��d��#9g,OΔ55�3�	;�j5�vmPa~����!���e�-�~l5���D �>6�r i��i���wY>y���ɍ�$��4S6�V�3i�&/I~��AT�_o=5�����1s��]����<��\�F;֖�V��ӵ��v��#7Ss����ZͲ����<Q��5XRUc���pRah�����T� ��KVI�]���'Y����U��+--r~�;t�}��' ΐ]ˊּ��f:���vQ�GWpskc�l֑���������h���/��$LH�C=� }a����Vg�⟕";��N�����J�z��UF&;{�DQY7�'���vЪ����YoƎ;%���[/���j�{\>}��¤�y�M`Ż�]<�"��**��03��ʚs �9ɕ����~�����(~��H7�LYƤ�a���G7ɽV>A���-��56U�K�Y�;��O~$�����d��c��y�'��0)�5�������z\jHr2%K���&?Q��wؽ��%�.�cN���~��s�ϐB�¹sPRWW_)�?�C�M-�z�����TGm��^욐�X�aŭc�F�(Z��O}xc�9����7h�Է��(���F�%��{y�����I�3߰��+l��]��Xܰ�+F���)����)`�Q�<hI��������Ia�S(�D6�c}Jl���O�I^�����1e��y�G?\]_��D�Tx�v�ȫ�Vѐq��>�N���C���mv�y��q�-���Y\BteU���^�=�L�{8�h|A����[�W�ݾ1����)H���r�m�NVr>%��Q�Chu�K�'�7�h~ˆ$�I��e���l���SD	I�Zs[Օ��ދDF%U]4=p/���	!yj�T�_��N��X���V5d�;��k2&	=<F��!����e\���>����z�$B�s&yL���P�$d�o"�K��%�-��D�a���p4�����''6�[�(>�W� /����m��7�_@��o V�R��>��Խ�,�2�9obleQEiU>)����qu�"0)�<��hΞ-�Č5N����V�Y�-ɟ��"&qtt,��|=���X�����-,�{1�����N�A�5��I�|���n]ƇD3;|Y��ޤ��Kᵚ-�ӷ�!�[���y��ɡ,s��	$m+QR)���i`K� c�:E�l�yuU�g���s��C:���R�3�=m!�r����ҥ�oS=�H. �N?�����_�%C��.�|u�:t�H����JD[],����r�z}�J��m{\�ޗ����lU,�m�h� �b)
���h�ؒ���L`lB
���W[GS.Δ�vB���m�<�����|v^��w�R�����֮۝��Yb+ ꀭ������*+SAN��Gb���z����f�V�M� v|�����*sj�Ȅ#mLJ�'�_>;/�KH���� ��_��:p�v� �R�xZ��6��Q�kL�f#I�3P�l���3?�qDޞAVJ5&�g�5b�����Bщ�]����c�aׇ�>��G��%���#	��Y���r�S)-kCp?�ra�ЖE�w5!u����C��y�C��|�5��71Ye#��=y��90�]��rk<:6��d�޼�QQQ��0̖Z��D�`�dH ߛ`<�;:򁚺a��H�]�j�W�ym�>zY��~�}$A��%�\�c�tDMj�\�*�oX��2f=V��tcE�ҘW��d�u�LF	,9�Y�@%SP��!ί�� �=��A��QP���[(�v��p|���R�m/��XN�")��`�+KN�j� <O�'�G�?�SSS?�Vh�6�j6#4�-��l7���C����hpQ��L��L����:�#��;�W�<�&x1��������ؘ��b<����3��z�zu�4Xe;n�m�Q�Ҵ�Ԩ����q���g��lN���t������1<����s��v3޵��-r���5�1���U/���D�D�!�,͸<˷��ɳݶF%Uվ.y&ʀoo����_1�ð~[M�����z�6���A��C�J���w7�ᱳ��~I�=���D�����!a���`�X�eP��Ю���z��tp���ſ��m�@��lQ�t��w���tw2���G͍��d{���p�H���5�H_o��uI��������~��qd�g�Z�\��N79�b���?��Qӌ1���ɔj�Z��2/�I�:�B�VE`
#���Ȯ��芰���]����b����Xma�U�گ	��~���e��	s�%�9�=��^�LT���}{5v	@kҾ弘�<K��<d)i�w�Z��~��2�떠�0EE.�k/�<(�Y'���2&1���w���eip8��k~�uz�DЌ����q��6���7�{X�5w��������=�`7+��"�;�K�F�;(�����!�׌�|/O��G��KR����-{�$�A����n/sɬ7 �T}��0S���,�;��h��rhx\x����[4J�D�糀
��R����j��g��k���F|��.�02��M����7���X�!��(˟_!m*������V���[��7����EN��0�}F��ӓ�v�z���vm/S�M�
`é��P����̯G�X�MfU}�苠�0���\�\~y�`k=#H�y��P�\�:��\aL�J��@�~�jȢ�\���^&��I��/ (�E.~���/����g���EU �z��A��\�(o�Ջe�iLo~C�bi�qq���d�f�H�E���Z�_~.U�!	�&���e>�2�@�_ױ�~��t�_au�	.�BE�N_��e�P���ey�;�6���|���8��'�`c�j�v����3�m��\�[e%[v:�D�M�5~8���X��~:�˙�ͦ�ذ��k���ډ��0��J����^�k�{���J{j�>�3w>:�|�9|��]F�ϭSE�'H��Ϥ;18Ȕ���o���X�ҹ�J��j��[�i�1�F�;31?��x��Gj��	qM����> ��v<8ތ:�A�b);��xq���ص/�5_*��>��&�����A�r1����[X4A���SV7ç�-�ȳ�Ê�N��6�������0F�N���'���Y*��*ZOX�F���7��Ⱥ�xV�����XK��xK]�{��z3+�P���{���Иl��Se0������!�� ��h�z��^x��4:�Iؠ�W��F������K��T/]��^��;.�i��}�"�'+�[E�1=UbS���ff�DF����IO�WUW7~y�լ6��͢�/�d��`;�[��Ubu[��]����JF~oII��D��[��w~�}���$~6�a`�������p����Ȃ��TP�3��s6Fntb]it��mѕ+?W'�O�q��d�w#��v�P��fD��5��V���U�jQ��Fb�Awe�����ȉ5��aY���Ԗ�x�\�M���,7Ϸ9���B]�O_�1�I�)������/���)��B-��������q���ME���~~0��D7�U��b ��gs{n_a�0���7u������-�%��t�ѳ��~�Qe��e��Df�aڻ!j��M��t�M�դ�̛!����[SS��XaTc��6�95H�]�E��;
���ȡ��e�����'�W��ĉ�����.�= m6^80G\\x4rbFJX7�Ka��2��?�lB��g�;�����CF2��f6o�l 2��?������O��C��ͷ�,��R�͘%��t>g �9��W%�����-~8����h��Q��Ͼ���_��:����iz\��i�$�)+X�-9y؉��z!��E�jV��$y[l��-���S3�`�%�wU�Ԯɂ�a{�!X��oap�9��t�T�]���`מd�$2��v�0���聕��b~�`��c�P�k	C�̤.+p���}*D(�`ؚ��R(z��0��h���O�����gE��*�s�_�z�Q�I�k��9bh�း�������y+*s��̭Y�wyP��S�N�J�����r�޵�4�,�3�qo�����Y��d�C���Z{۰�S|��+��ilT�4�)�o��m�>�sa
���{����d����M꤬��N��{��\7�g� }ot?Z;��X�53!wC��4G\�<߭��,��~KԴ��v��<Q�Ê��au��J�斈*�^�v�J�\	F�0�f`d�8��=e�a:{��E!v>����p��)�G��ѡ�'��ÊF��_X�޺�¨�v�@e T�)a�p]���	�!�ޘ�$�N���(ퟦ��J��wW�a=s�pQ..�_��hE�m$M
l��w���m��e�(Vo��S:�"��A�}KR��~��vq��t9.�31n�Dg&��X�p=Qà�����9r�щF�d3�IJ�k�Y�A�����'�G�!"��$�UX+��_����0-���:9�!ÙuQ.(�̺O��Q������t�UϪ�r�հ�a�7���/��d�4�>i��Ɛƭ�|ñ#��r�-��|<��ܦ�?_�>��]\�V�U�֎�+o�7��Џl&돨����V��|��R 4R�7���
��mA_P	�k���'��ǒ�N(1B'��.S!ɜ��؛����v��.��{�@�של�o�ݬJ�����'���%-�<k>DvAz��ZW������Emdј�����_7s�}�`.��O`��D��=g���0^����enZ�1T��RO|�R�������O�-����w��Z�^^���h $��P�`�0�#�`u�F~��>�)XIq���ѳ�W�\�Ez=9���}�Y�D��p��x����P����
�4b�z�Ί��><,�k%�xW(ˏ�+#n��= ��y�
{�N�|�}m�vBx0�j��3/��:���hxt�X�~;�	�&3�>s�_��7wh*(|��5��r\;c��;XS���YU���۠���Ki�HA��Ֆ�A�h�d,�
�Ǚⷂ����voW��""Bn�xbg=p\Z��
�[JJ
!��G|�aK���}�Uu�qy4]Hz_��x�TC!Y[oD�j.j�l���qz�Opy>^3�>P�b	X:�p����cll�JO��U\(ߋLKx��<մ���S4rn4555tfePB�*/��z���I(я��_�k,X��[?&ϗ�q��&a̫�ZM��w��P7��d�Օq�Ё��Ns�����;+�'��s�kk�OWjgϲ�������^Ū��9��T_�^k����jB�����p�<���[��܌a��ϟo_S5M-,�xx^��gZ	�g�+��\?Zݔ�=�!��{�/�oG�i��~B0&bc+J@�uu?�spL՟�w�׻�����C��~o��@���:��������u�j���Cs����#ŔC�AT~gg'��[+���y(��ƾKNM%�ۼ�HZZ:�ס���3:>[��ׯ6I�	II�;N�,gO�o^O���ޜV�Y�A8W.�VY�+�ܛj���R(������deŁ���p]��dU��]�G�$�F`�t��p�Bs�����k�7��J���\t��q��q�j�C�(k�E��m��3Z^���ˋ��R��!e�%�!hi�n-�y��Ã^x�f�U�p�И�ZB��QE���5�p ��bs��b������w�!x���z�� �db�0|���,���u��D�E�4ld'hi+���k������������mfq���:,�o�^��3��
<"s�yX����/1 ��ǐ�[��y5�P��*��bM��!�XF���9�����
*��Z8��Fip6�6�5��tMm���h��!͵e �G��|��e�!�]�)!�{�E�з�8Yi#fo_�l-�.���~6��G���z#� b�ye�DDN��_�{���_��>�8�zK�,�_��FH�����ɇ\���gV�|EG��<�1���Q	)��H�������v�ɿL�T����e���
���OG�TF*>?�g����=�u�^�+g�{��#����Ys^iRÈ��B����K�Ķ4��BeO}�4�a���y���n,��S����_!Q��
J����B���K:M�f�����]}V� �����.���kk�qg�͵�O;���D����
�4�]A@ HP�Hҫ� RC��(�{G�A��A�� -t��J w�����s����ݜ���}�=�<3����Бk��Ln�Zp=�.旐�/9�oڟ���ƶV����"���2�=��$ߧrNq�9���2w�|w��ר����T��&Ӷ��MR�G7g�{,���gl��W1�X���_%z�"�����-9�`����_^ِkf��;/�s���9B�^i2�,��&�m.��hN
y��2��ry��/��ƫb�L�����o�V.��ug5�"��x�y�m��N��'�)�)���-������az�H��}��Q�Ļr���3Z��̱�g0{��	��*�V�/�u*v�����1�|{�l1��.j�ɠ�.�[�1E��æ���(���$-����=ط����k,4i�||`��3Qi��s����師��B�S�Er&Q��d}rN��	���f@�g���@)[=�?�2�ݿ�&*���+�}��Y\\,"*��j-q��n�%&Ջt`-^��o��W ���7V��ƪ������۾�HZLѰ����B����QO����Se2��><�����h����&���������S��ތ5��Q��P���-�LHi�Q�]ޗ�WA&�3Q��Hr�U([+��<մeҷ����$;�k���X�ys�a�� �b�c�.-�Lh~tݟ�t��)y����]ccc7��c��5������F�P[����~T,k�:�mu�t������[y�|�O�l���]�*�/�b�$�(��Oi�`���q��'^�e��D�-��$�q���Qjt;����`�	�G�؇���s��8H�3aTI?q����`�39�����RBɝ�L�������x��l)���*k�V���ې�O�W��L�e��8�s�K�ɫ���@�S���-(���ȃ�h���O�e$ě%?u�1a��Sv�m�cwĚ��La��X�ZkV���s�p��T��93�::����w���'�m�ȴ�4�������kWW�t���t��'~k#��=��l�cv5���ו��MT���"Sp
QśUo���a��'1�O�=����{Qk���
����7��Y�zEE�~�7a��B�aޑ![gG̈́~Y\���pe,�d��w=F�+m9�l�Oj�3����4X�mxL9�	c�������r�^
��_
���.'�Z��8��������C]{�1�<���7�D������)�Ϋw4����d�,�f�/���씙���H�Iv:.����˟��Lyeanp�⹫���y��+���1�	��je�\}�bO]����g+��Q�Q������5u��b��d��=ςPp+|=v�;S�C9U}��TX�5ex�*kc�~S6Y������W}=��ӭ.eZ���&y�sx�0r���L:�/�(H��U�^+�-�t�h�Vii�?4��(K��>c��(W�����8�ZA:eE����-*.E���3�[�M�z�uk6��d=5��]w��xP{������|�P(�w�t��5twT@�����M9��n���&cuF���ju�Y��0�k�rnM���S>!-��;DF�.˺n��ڻ{�;�5�#����{�u'���S�j�����t"A)L�;��G@�t` ���hű��o���b)��Z��jas�����R�<���5Nt]M�c�y?N���d��2��a+��Ɉ�)�|+��)���ͩ��.���\��lD�Z�[�����'Jy�o�Ve�[[�U}Bm.ȮU��g�^�3�)�f�׈��,����������!�x��ֵ�Ͼ���1��l���P��lױ;>�٩@O�˯'/'.�S7s;%U��1�P��^��c�vD�񭣘��C�˃M�������]�k�,u�o
;aC.J��~<���zÕ���������h� .���(��,ش(zU;`�3J�ZI�U���e�ƴ���{�Q�ՐLk|+A{�C���k��h$=��p������@5��{�p�U�1Z^_�'����KH�k�^teY\�u��P���i�+��g�h�^G���UCT�J��/�k��y)��6�E�'<R�za	��������]T�|Rq�����1o�֑Z��Z��-���%e[)p��#"(����JJ�`�7�u����8F��hx�}{�Z��)9^�"}h�6>�$!+mo�Y8g��l9'&6��\�o,�H��6f�,<ג2S��=�7��!(��������b�T4t�p���޿�O�+y��gf�SU�2U)-�!�NҾF-%�{��2���w����U ��*��H���Zt�|o__�f�'�`ȳݰ�^�������ԴTۣR�m5#7���z�0c��E�8׳�5�ظB~���z\�b!�c�֙a�l�ܖu-6duoxh��d������}G�=7�5E���qs�=ѽ����$7���K������)��/1�,3{e���+�,IIIrb#�m�'%�������i���ui�[;/�Bo����`���ǿ�"�&��f�}��
V��]Z�^8��9|.�sĘ�ƾ�q������m��r��˨��g3���O�v�gEEE��KŚɥ��7=>�W��-J�Fvp<���4q��m�e�\�<:�����A����M>>��s?r���g�E������k��u���Wűz��L�����(��:vj�j��f}@ژ�ԝ�^�E��	:�כ�%&}��!�UUؒ-�ћz���������	�E�O���y�2�F�W�����~ȶؤK]437	����܉�8ڙa�a��p&RD������s«��r�e��1�e������	���Q�<�f*�^�$�S��RRپ>>\����/�/��T�j��+!�|�"����#*-(t�ǚ'��#L#�kx��ƒzx��E�l���z�o�"t�L0��x�gD�&�X#"�jVPPд%$�(�������r��֝�bQAal���/���B�_�6��YT�� ���@��+��
%�1Xz�Cj<׎�Q��R�1� I�e˼�F#�<F�Tvo��f�ƅ_��|���2�-�[C���:E�ׁ����{e�+'��-!�Zl����u���>D�3���P���>]/ 8?�u��7zЇBB��s)�*-!v����i�^:���MuJ{Y���]�"�����x~�4�Т��R'�R~9� ���{Ff�ERR��������?�l�I~}�޼��4�B�*9[�0V�z�U�/�<'�\~���,�R
V.N�|���W�R���ba$S.�|����S�._߲�ކ�s]3��w'+�+�����<h-�4��|��.��gW'��q�7�s�?�p�|4���]��*���2Շ�_K�f��Z���z��h�s뱝ݻ#B�㹕p���l��������1Ny/0G�Z�Nf-�+I��sj,��¥Ug�d�J�l?G�.����,?�wEi)PD�I��ܹ
��mw�v|Qt�y���s7/��0��}���N��«V���弪L\�nf.������o8�Ǔ3Sw�ϫaO������W���mgvTU{���vJ��/���Q�S�Ҫ�2��-_3W[�b����w��V���hu�x�hXr?5"�8pg.��[���e y*������\1�/�4��k%�/#��⾩��}��GĹ�L"��><�]������+��e� �i@
���:���b*��ꇨ���Gbn���(�A6Y��i|�bv���u����A\כ�����*&E���+�q�o��?��r�70h�K<Zl"�GW�KQ�oQ�:C��*Vڟ�1�l{ܰK�.�?#p1ƽɜt>�~�Х��N�&�m�ƮYK�c9'�}a�x�k�A�^'�����~�������.������*Hdff6��qRڇ�y��֛�`�	::��i�Z��m]���X��j����5��0k	��h��L�S�+3�K���n^`��L�7�t���A%l@k�k��V�n��OgZmA�C���l�Z�(�����ȕ�yߕ���α����C>��|����Ze���9�Sq�(��˩���k��P�R^����n��p�@Ս5���KUؙ���>9M���[[�����+@�I_�����w����0\�s��HW������G��G���kp� �'�ؿM^�h������H ����uʝkq�{"�56��$:KMW	]����!a�Ȇ��_G9,�������b�A��X-��=]]k����t���x{ץk�G�a�M�;��G���U�HO�����fC!���C3iǅ���xxy�^���m�A��ee�4M���Ȟ�nd4�m@~eP>h&���t���{K4��>�/t(?��ܽ>H�Lܛ�{}�`�Lf��뛎�<)lt���n��I���z\ߘn&R� ��ܡQ���{�@�b �|��÷�Rls��V]�����f4���
��T	���*���*vZJ��xLCN+|���o)�91��62� űKo�c�K8����W�����F�a�A�m�Ɇ[R�4�(휗+}2� �*��M^+��n9<˯��Vڗq�%_��y�uq݈K/F k�D�C֋����}%�xȒ���o���eGgqX��B���W����y��Oţ/�Z�g �އl��K@�&Ox������xT^ʗ+8^��������s��zc���X6�%���P�Z�	��Ǘ�\����@H?��g��\H��\��s���L������_by�����g��t-1R(Y����R�4�m�y;��8���㸼�V�����r=�v��TO)=���6�X��\��*x8���n�cd{�۸�O����9S�4��@!7H�MG����i>{�\vM���]���u�ܶ9�5E��jk{{��JN���Ae��)�fq�Z�x��[B	le���۸�IN=�+V��x!�CA�*ЦJ�w�{�6�s�w7�-��ͬ|�%	�VLMq��4�(j��U�1�95;�ۈtť��+C��E�'���/7���Y�y%�Z3n�c���:��
9���ٳ�T�j�q�h����}���r�ͣ�!1��d�����Z���8�?���%�4All[���
�=6�����W�8�}<��4��Y�φ��s�;2�یL򳒲��P���ɺi�_�.�3&~�g���>���4a�	��_΍�\����<�'%%e6ό07��ݽ1]8Z�O�T�`V��ds��Ƿ/�)����/(Z#�e�	�x1�����c�N��r�Of� vP&�&Y���r-�_y�Ʊ؄	*X5Fڰ���|D�$O?�΄0��b+%%�����R]Ĵ]�3�h�ƈU��I0#��{ǘ+������݄���o�Ĕ��l��M"i����ʼ�X����n��:H!(��|׸�B�a�Uj����&����N����[����AK4�\�f�_�#����S����;|��w)���+5�;2�<)��Zj�>����\8�F���������KVψ�
�N�*!]f��g�V8L��Vm�z�&�$N��Qg�-�A	)9���dN�Q�-�>	��S��g^�/[�r�sȋ���8��l7)�!�^|��� [��$�y.�CU�~��}�V|�Q@��!��xГ*�|g�ۂy�ש�~6daA�H(;ؕ3��W�Yf��+7;y.,�Ը82�S�>�z#_0ao���'�N�V�?PXd�&�S�;x9��i����m����m�HI��}�Q�_JI9@�+[��/bS鱕���O�KY�|0|n���W:�]ٵ&<L�����[#E-��3��ɋ��J�s�"�Bl�GӍ�_�����>�)�=��� �Ƙ����r�k�#Oó�KVX�B��.����>��I	�����X NQ����b
����
���ι�g��'��pn�.E��,���u�����-�ԍ6�]ʲ͆��/���Tn7ݑ�w�t�L����r_&������Sz4SR�ϟ��;:~����B����GS��S�z��?��oI4�m-�QLwA P�������*>��`Q���~ 
v��0�E��0�B�J(:��}󿛬����{�,��W�ڳ���0Y���p�������>��	tC򆤸����ԃR`i)���5II���AOP���������D������E 9�c �	���99�:�A
�f/����l�y�tt7U�=r���yz�����9ہ��X�����KJ~_�JdD�20{{���W�����o�玗��#������I)9�6� ���8���>0/89IU����� }����&��4�tU�Tl#�PK   �p�XT��_�  K�  /   images/aa07afbd-658f-44ac-9cd7-fcb1529195ab.png 1@ο�PNG

   IHDR   �  �   �$   gAMA  ���a   	pHYs  �  ��o�d  ��IDATx���%Yvv����ʴ�3=~v����X��p\��II�E(B�w�I���/P� 1DB4 `�Y`ͬ�===��?��^��1i^U�T�T�,�կ�|�7�=���9'w??~~|N�ω����v���~~|n�ω����v��_Ji����Q��O�������߳c�>��]}=����=��ۿ��5�1<�����˯��qЍ�����ko����#�A��?�~��-j����3I|�=�vnynoou�'�����+�^�2�m��cZ�<51O�eXS�Mz�-@��E��KM������S�������H���G)���ަ�$zu)�+���ӻ	w����E��ۙ�Wh�)�SN#
t
m�籅��-D�Ə1����c�2���ϣ@��(�)<�>���l2�*z�U]ǅk��~��;aT<������إy�����3E|��w.5��{o�M��T_�M�A�E�4n\S�i�����F�X6>�^��jʔ��t��[�|���kz�3�%&V���:�Z?�x�>-#��п��`.�kǝ��t�ϰYj"<�1�h�y��\�Y���lte�f��*���Ě�bI���*;Y�T�_,���>��G�޼��}�����?�G�6��w������Z��?$���6q;�M\��2&��,�9���_̃T�W�M���/��7�.D<�i_w)OR�7�>���}�`Jx��vJN�JM�� �~yT��o,���j�����������;w��:>w�#}n�o4��G��I�{���9|z�GN<��/f�.TX��R�_��Ny��v�$?$� ����'���wm��O�A�4$��;�
�	�4�Eu�XH�q��!��Ys���Z��zp��?�����������v�[nY�3�[�.���dޟ̫�9����8�OIu�x��1�x�ӌ+�.;v]����`N�v�`&��r�~~?6͹�X��߿��^�z�g� ?7�K�����՛eU�/uS�1)X7�3�&�&t��������o~�1�αM�r0�(�q~�:�~M&����k�a���_�;�7�~\���"��T�i���裏�Ս7����\��&������U��c�I�us�����ɯO�O�Γ�)����)��a�J~?~�>���)���K��h����Cmi����%�6��%�6�����+W�����\�oww��*�I��^ L0O2�0���~��lW'�p����X׉"��Z��^'d��}UW��ul�� ����J����)?�$�n�E���?/�k�h� ��p�Ţ����c��w>OW�gN|������_����Pxތ�b��q�pX��a�1�
�I��G1E����������'��g'�K�Tw��>kߋ��5:Vھ��Q�|��4�7��s������t|��q����W���	��[4-[�4'_{��[[���kD��3�_����&��ծ�穎ŋ�O�Pv�V�H�u����i���v��R�o�(���\B����e��S��Z��~�-�}��ݝ�7o���p|��G��ժZ�.M��h�΃�bM?�L�Yx�0�����$�dz��$K��^�k�}����j�;�i���}B��%�'������!�^��v���>�2"8?���i�S3�����r�ٹs?�S�>��3#>���Ç��HM�M��F"�kʒ'��@6�Qtaс�abNOWkR�hz��Ε�!�0$�l4r�X1�"�u��06_hjG� b4>�i���YyD1@x)�����U��T�~�1��‛�C���Q�sÍ)�ۼ���l�V� "�9J�Z�_o�e�cS��j����q���C������]�u��4�o�<5�-t�,�Kb�5���$��÷�q(��X�X���aDBj"ܺi�@0݃�MVMlvR�i<$Bۡ�&�I$>��_��y��u�޿H�msD�bN}�)	����m�'�lM��GtN��$�;�}���d���\���������g||&�����ǯU��eX`M]���x��ǝ��w�K^�#�3��2��])��)q�:��(')[���5�"���7��_���ɴ������q�j��݈��zcU5����u�|=6�/�}n�m�
��HֺpT!���4.�D`\��^|��fI�%(���r�t�^�~�p���H%�{�ҥ}��	����^MM�M��/��1��!�%���]��5�n+������Ȗ�v��R`���Q�3��sr��NU��!�~4�N�EV��t:-���=~���<���cz�.]������><�����𷖫���*}v���`l_���0b�Y�s�� ;��PW�_���MA�Z�W���lL��Co��E|dMW_�F���+��k�ԭlHhk.���_T7�u���k<8��+��Y�[t��HG�K��G"�~������w���A��Z������n�����b�G4"����u��Ms�:am�Q�����#�ч䘡џG#�nñ������� �>_�JL�����w�gt<w�Ͳ�H��%��1�+�J���N򇵿���� **��	��n�W����g�T�;�/�[�ۥK�������^����g���j���ߤg��l�wCW��w[����:�:n� ���zF�]M��rY��r��w���2������_'M���Gu=�x�|��k"�'u�i�NL���A���p�q]���4�p "�E��;綶�����ާ�}^����λ�}?��|qtx�6�o�!�Bul�v��k�*t�T��ڧW�b�A�����"��\�CnQ=�N3qn������vw������?|��Gj~�&�4�����灈t"F�G�k��~�\��OR��u��(8b�:�|����/���3
�_x���۷o�]���EY�7�6�0�kE+CϿn��}��^�l�y��ۿ�`3��&SLbSU���o��o�ψ�=7�{����|�+������RW��W%[r�Ím�1�G8�T�0���Ё0ݶ���+e]Y7�k�@�D���b�����]9�'�^|�㳜�_|�����	U��4�+d]o�,�����<�7����gO���_�����q�n4���r�F�)>�P��>_��$ݿ����~ϓ��"��H�~�t�l����v�P)>a{��]=|c�Y��O��gM���yoc���ln^xןq�w����X��-��8Ji���Ct\�q��sO$.{�'}.ĺf��{��֓��O�=��j��ͽ����I|;;;��z�Wǯ51�7�J�ԝ�֊Ǭ-����6���w�tAS�Y���Qm�]�/��8(����\>�gĥ��p��B�p5�5q��uQ�2�=W_�2�ț���a����������#�jN�#��U��-���m���?��Ӕ����W��9υ��"�Z.�7i�^6�cǩER7)8�j]���"�O����[�놜/A C�DᏳ��s1`�{���UUU��������q��{ظO�x'�uI ���ߘg�ԣ�_|w�{��m��3'>@����WSl~�&y{��8��l��@)��z@}��;Nlv��b6v�zT2�NiU䣇��t��NG�$�H�Ś���64"�zu�nH�����18�ܳ��oZ!Lq��kP����t���~�q���t�����9gJ|��a��keY�C�M/��>F|'�8�pP{�'�o0ɡ���c��Ō���m�<��%�=�c3�y�B&Z$�����#�!��}�c+��sN���Y��op�&�լ�_������7v�m��Nz�=��L�o>�_[������뺚Ş���Ҩ��F�,_׷fmg������c����M|\[�:O���˧��38���ʱ��¢���]��T�͎|M�6*p]T���3�7g�/Bܻ�D�U�ފ������%�~����wf�G4:8x�jS����v�UJxՇn#CL����V,�9Z��n�{�rݗ�;�_q_p�|T��'?�F,�=��#�A�N��sNyݴ:��O.������	�F��_k�}Rt��i^7�����z�x���{Ǚ���� E��~!s~� �E)�\B*L��J	%��ۋL�OR��;���YkɐĽ�HR.�;�?gr=пh�����Ń�j�㱿8�)�l�&����m����ΦFsy��!��[Pl#]�O0Hl�Z�j�镸�5E��<���_]6�7�Ų���ݣ�n�~�o���w&�G=��{��XD3��6��e��7��t+� � �����=M��E:dUo�}\���=�IF��9E/3��EH��Խ��3�๸Zp4��m�K$rs��VH:�p��t"g��}+���;w2GԳN�z�q���Ċ��*@���$؛����u���gB| �V��7SU15�HD^����]��2����"�ѷR��_�����+9
�{+�5��G��&'��2p�gU��[�|�>����^�O{�u��y��o�s�B��ʺ�Ta�!�����	�|&s��3)��K�hM6ZH�ꎩO�z̃�ۍ��!nT����Z,��`z�g�����s=>5���?~�Fݔ�G�y�����r��?<Lq���|憑@Zh�z�-�O|!r
���rAFu`�iLｶ��������=�z&�yu���̇�06��af��s�nB��?�����t�skܴ���t�����7�M717�3<>5���o���۴�_�q������z�I�+N����D��RN&��`P���oI�}-M	*�Y`B,������S[>��Ŭ�;Ғ���g�jXɾ�<Z����GI��=K�����~��j�w&��6�p4?�zV>�t�0�W����zM���ܙ~�ݻg����6�r��ֽ	���{��"�������O�߿��,s=>�ts��"��4�k��Ǝ㹞�C�1�����m���������z����8Y����\lL,��/�_�0~{:��g�Ν�����O��~kT@%�Ks�-�+wL�b~��6}�U�������L���͝`q�3�j��+�G�oL6&?�tFS���������oC1%]/7�O�՜�X���0A����g��$"���~f�D��b��3g����N����4�Sb��GS��i^j��>�>xtp�џlm}zX�����࣏��.˿�g�Ŧ*[�&se\nM-�1�w=u�k�ר����q���M�O����X� ��ܹi.��ߘo���X.^������������������x�od`2��Oq~b���$��,Pt'h�;?��qo"�w�����~&1�/��>�g�{�����_onn���۷o�����?<���t痳"��bj�d��Uu>i~���1��A�ωY�Z�B��.i��5�O�׍QT������w67���~��G�s�8�6U�f�\ϫe[id��J�>�۝r�7�u�Zw)tn��w�\-|=������5(��`�=+�-w5� +7"ݯQ4�(/h��ͺ�u���������}�gn�y���{:� �hs��{����yt��?����f�r�"1���<ط`Yp�>G;��#ٌ����"�=�kI�����Ȳ�'{�m����
����˲�����o�a�p{{�����OE|�L5��o7M���M�F���Фk~m��u�s��uC��`Gz1N2��:KS���ܡE�6cL-\��<ި	�&z���:��W��.ӳ|u2;�7�������77���S�y2v�����{����꣏�~����:88�ü/6)��"j�W]n��JG��s�>+�7��y�%���*]f@w���>��E�ln�����Wb"�0�[7�B]��\.�Ay��]�S�1~*�����|�(5�U,��k��8����\Ċ���j��v�5�'�&e�A#��`��w�TP_�luYh��פm�WG,����ܧ������b5�>O�q8���d<�����O����;��g1TU*��?�Q��W���ˇ��������~�6�E 4����\�H#7$�r�����I��D(B]�Pa�Z��g����C�7p�:7�s�#@;���dL���������>��?U��g&>�&q�W���2�y��~�����h�b7����Ƿ	n9�n^5�#�UK��[|!븪����"�s���\F艚�jua݅����w��ܽ�h����Q��$�����m5M:GD����(�<����)h@�L^P�\�&R�u�z�7*�����;���[�'�}�ap,v�{.��,�%(HQ���{}Y�~�h6{[��O�x~f�[����J���%ʛ:���c���k���])Jf�S]Ŋ�����A�œT�Ib,H!�,�b.�P�p?�"+L9!-~��{/�8��
G��fRmJ����Xp� \,H_�b�ج���${�&~�`��$�%�,<�4@�xթ��2��B�������T��2�6`�H[�(����ZK���Z��%�����I`��lD�yL[���kE^���x|���c�S�D|4�����[�	~qJ���ʜ	���3?����]���5(��5` �����r=��¢�Ɉ��rŁ�������颗Bĉ��2!j[Lm�����@�����l\~�&'���ҙU%1�0Vp؆�ԌH�4^��H�(W+7.rd�u����p5��.(��P��៰F'r§�iL�?��T����C0j��������������{d|���S�ğ�������k�د�`��(DFŏ:�Q�W��"��,YZ-4u�D'a��u��0��F|\j�,�y�"n�h�z&��a,�C��vqh��d6u�[�����eн�p���r�h9L��	���E)�"�Z��xc�mn�\1;��pfI��{U.���t�#�֘�o���r�k�_ǳtA�y2��s�d��ug���qf��7l��˚�q�#��7/�E]Uo,�����s���6��̑�g"��L�IO�5��K"2�5Y�yOl�[K�� �Uf $+���ߴg��P���j��N�GZĲ����b
��R��┓�[����S?s��ҥK|�&u�=��J�O[,�0�����u�0s�pT�9�Ͳ-����ϟc5�]N�l
l�|,��<փ�=��D���2ݐ9B"׍P4�t1���s�x�l�WU�)�9�U���v�36�Pߒgc�Q�B�e�v��/�����X.s�Z��6�]����<5�z����͘�WB�%|:�MB�&�D�+����&Ca��>��ҝ�oN������vP�®gJu`�X�пz����"n3q'����b	Ը�7n�)=�~/ž��%'��I!n��b����k7����,rKT��%?�s�:Ys��ٸp��{�75��`�k��C1�ʸ��D��dJD��.^t#�>bҐ=��̩�T�\dS;���5��|�� �H��1��w�D/|�n�գ��Ho}�ރ��L��S�����7{o�,��Z�i��`;�5��W�����+��S�eRj�FA��)&c&�բv��bI�Bu���>Y1b�l<%Sd,�X|y�%���(��d�,��MpWDV�X<[��c�O���	#"�UŁz��ZF���c�X�@��N�F����xg[�t�)[�rA�Sg�ۜ��6�Ѓ����L�/|n��U�J�k�띶��[UU�}��o��w�>�O:NM|$>f4/�M6�h�ٚam�6du�*�t����߆��l��Ik;���DHZ�E��>��| 8v�dāp���vy1�7�qx� "y1Hp�V��K��J�tj�Z��BD+��x2c�*UH3��A��J��ܰ8Ŧ'\-n~H:i�b�W��C����#�i��M�d3q��5ǥ���FθTj��K�p}�[1%��ahζ!��S�1���W�w#n�O�+����Ss�SM�F]��>�#c��}}��n��$}�����'�p-��)�W�B�����9�ʙg�$}(O5����� �E��h�=Lln��Y��rp�-�«ʕ:|��oEo��T�q8�Qe
T�t�u���Lgq ۗ�R��
��\O�q_�|�Ѧ��L,B'��ZnԉϞTY���I�هuf!�1 ��}�$�5Wi�~�t�����6yj���,�$=/��?�H!����<k�;���?L�d>(��O=C�3�DXDܣ�#�W�.hd7���	��?��#ΈP�g�Īk�)b�����e"��d�K�ש�:1��/��L� JT`h^-�7��p�<Q��g��suM�<��{�?�;G����l|27�U��4ĩ		9˹B���Hܢ?�up1��8����b��� ˫�֯/��v^pC�~��1Ϻ��@��Úu|M(�	��T��H�$�*�ml�`�-k��JO��FP����Q�o5j�;�/~��HW�QPƮ�)΍k�}�Z�Q��z���c��d�  ^\�8F2��mz�
v���uD���?�#(��O|����.����羭�B< �,ʋ-gG|8���	����
�OB^�@�RO`p)��@�Yf��D2'���'~��&pB��gE�G)C�D-��t��8 Bk�*)��C�ki���Y [�5��`l�"�Gy`}��\wF��*����L�(늸�����wըs�Ĥ�1r��5�d��������ݭ�����>������S���Mh,WIO�)��_�4e�D�J�X���g&����'�������I��'v�H���p�f�$�"YYt'IةS'v��n&Nh#x�	OꀉѢ%����ɸJ�`�UD�ә�#���M�muN�B@�x�pVKm��"��Y����S�vѴpY�������''��ԕ�~��uxbP���F�;NM|t�Q�%�W`�]�w�_�l�~�ayصl}������bp(p��I$cggǥ��m�Ƭ�-�K7��t+�tGs2DhC��F�0�Q��3�E�lwF+�j�G�n\d�K��AFH�V$zq.�=���L@`,Ʌ3���ə8�W�r�uv�9�?��W����X�Q1qK��IeX����[2�g^�U%h:D�Ɗeӻv]d��L���ܬ��$U}ݫQǁ��$c��j}�qZ�C��W�'Yz<mw����=aG�NT�o׷���*�V�_��{?fݼ�$�Q6��9��K��da̶y�8��G���i� =��N�����C���G�upbmR��*I4��p/)a�'W��͗w��m�?ě�	R�>~���>Be/�W}ú��Ɩ[���ZSw��7�O9�ZWW�	]�����P��s�u��i�k� �(�'�8��Y8�$a�=����N��Ϛ�w��<Ⱥ�6�֯�ǯ�3�N��t�1N|w�X��[��(cq��#W�+F.��Nc2�����p`�l\��n�pI��d�|�����y"-�4g��q�
�%��=�aG�sď�I�Ūd�e��J�/-���5r���9���a�F�'̻O4ޞt��	����u9�:�������%>O�,�cEO�'׺_�����$=��/|�;�a�(�Lfn:� �n#����ʜDnFę��\V/�b�r[�q#('2ߡ�d����!ȮzdUEW��$���p��zO�R��.�(~�Z�� �"�9��t�V�C��FN�]Țl�f�ՠ�qe����Q��Ӑ�|�dN���3�ށv#�9q>�A���֙���x<��$��~�!��w���u"�#�	*�ޒ8s&"��8�P~�s� I�,W��fL ⨎��käۿ��}Pk3r�mN׍9
by28A~���q�^ޏ=�R�|��\3d�.�+qf���3T�Ț��)iEWp	���Q�4q<�ad�#ڜ���y>#�!Ӱ����=��F:r�6�FJ��ppTJ�8ߺ���;�#���_��=��s\G�,����8�Ey�:Aw
��߽��=��wWo��-D�jY���%�F'�		�Q��xʮpP�,��@h�0LDs:q�2
�9*i{G��?������7_{ͽx�+H�c*�pH�'"���_��vǜ���I�U�?�>�ӏ��Ś�-H�9u��S=܈&�n��\9�ķ���q�x���#��k����'�8�d�A�A����X7"�ȅ�=�? ���{���MDw����ws�qiYt�$Q�I��u��}��b4f�	D(�C^¥��u.#x#'ә�?���~�T�w_��{���ŋ�cC=(��<a�.�V��0��m�5��D{��U��M�5�݈��B�1�E@�M�x�'>KW������?�-�L����a�+����j����.�şnm��|w�p��������݃���˯�B��rW��3����)
���T�He.$g�u���ge��z��c�L���Y�,�j⬤'^�r�M76�ݏ>f7\7_��?���ܶ ���9qM���Ij�gy�qX�4��Tǩ��s���Be��t77�A@������%��н��~���<��'A��h�7H!���+n1��3#��P�\������K����x�ݸ�����t�Z�e�>ы�r�U�D��M�/�WK��t���\�*����6YC�^�p��p��b�n.�F�ܹm���|���Cw�6IE��2=wΝ?��j�6�~nhAB�p�z�r:�y��B7�?���O<Z��e�}�މ��%>��P��|�����;�Y����o�G˦�\���Q����7���8�EO�-WG���ͷ~�-IB�}6�v׮�@:�����t�e���:�%#����W�W�_gN;*2�b	�=1�e��镫�YD2ƆE��\�K%�&�o����[o�%b���͈3_�{��A���Kƒı����)z[7�k���Y{w������N�j		�2u�=�ъi�i q}���Ϩiu�߭��H&dl QMQ-��/�a I6����EnX�P�9\%ζ6mPGh�b�9w�]{Sro�r��������)�R�c�qo_~A�t�J`΅��9�pקם{�u�6�k���e5�Z���n�ijA:�|u�OK}O>��ʧ">��j�"�9;{��^q^��7�{���0q�ˡ����z�[
ulD�*/<[�$W=~H��:��m�5g=�e,e�dqZ�J�]�i�.�qjeTw<Tbܾx���b7�HCo���p���:����SoN�)8��	ֲ�3w2s��7��/���O��Z��z�E�j���'�ly��N�P�e��軣��Z:,F!�$0�ឋɈ�_�a���f9��h�����8�/�mq��~���2���r��M1a"����o ��֜�i��9�*�T�ݦ���dt�'��3�*'�Wk.���|z]`�Z���yb��I�7_z�g�2З�L�]��A��Z���o1/�
A�I�_������qUV�ָ
p#�>_ci�b�c���nZ)�%q��-N�|�����s�d�����nqx�:+W͏�,n�K�A>d1�w��:��;��;󧱺�����pV��\?��?�Y��בk��쭾�1�b�s�#�e,TN�����&d"W\�����Վ?HQ�0-I:B���q���Z�҂��dޔ������4#N7��@xF�d�ǖ����ےNPجo�G7�:��Z�A���,h�O&�O)�}]zF
|�#+�eb/szƧ!_��U�a�����y���˒\���	C�qH,jiY|�5�n�Xuc[�_C�BȽ�]�W^"��>�^vB�6��6��� 	H@�1�y��t~Iτ'X�-P���u��N6�d6��3�N�_������\��j������!sќ���'��ǲ���7��ʻ
S��axN�<,OdpIs�gi$@��D�(����l��媃�J���^��ަ��������j7M�%�3gKA Y^<։�S(�<�g�I� �r	��YKC];�6��Xs��бx�e֟�~���I�Wib���E8���lVL���X�<�7F�㽟��R��zO;Wc�BUk�����L��愱�߅�뻊Y'�c� �)-��,�oVn��o�Ik���������O���<���1w����"��{�%���]���<C�Z���,B�Z�}b{����uԾK���3�_��!�������e>zs0Slu<�bm�\O�l��ec��+qx��b�2.%.�he�|�#�^9�޵S�s��d�G�{����\������զn�U�6������T�ϋ�;fI�u���a������c���%��?��#wb�,BY��$Cq�s���}�|��t�m�]���^�����0�K���]+�!��b��?�Ѫ!㺿�lq���G��χ1��~��~��������څ2����!t0���z�O�?	\6"����i���]%[��D��v fu�ƟHe+o��N��8�����t]�]�� b��s��U�T�(&I򉮫?s\�������7��̲h�d�U��s=�n8�v�dϩ筯�I�ѺN��]!!%b�He�9�qZ���*�'��������]#�7-��{�����N*D_�6��v���A�:��o�����?�u��#������s�{.����A�kH>)�i���97�]�%N6B�@�Gǻ��D0��띎N:֍���q'�����캨�w��Z@"b�yu/�0����D]�����z����9��/բ�gu��6H�F�l���-QdƊ����Uib��4dW綘�}���^��;��'��D1�z��d���>N{�I!M�J �sF�]W�[D對9&[6/��MU���*��؏]I����G]�c҃��q>�=�@��yp>0s�L��]\]��Џw�0P��7Qk�t!��k��$���{%��:XWڂ7W��S�H�kI=0�^Kx-GU����C�T��S׃~���'&��u�`��w�a�E�3�ZA�u��q;��{~�(D	�G�?���O�R���]��@%{^[�i�Z���r��\U(�>�9hk#�&�L}���X��A|4���w�o���C`��9�跶dQ:�߰�.W�QlK�umw����\�W�J:�\I&���_� �n6-�����œQ�"�wc�m@��J&�*�G;qժ&�+7Mm�G�\9�q�Is��< u�˥m[�`<�^���=���j�d�ǜǌӳ 5�~E�	��7��\�d[-�9b�O>�n�}!�̤眈����.�3�xh:�f�VҒn���}�zZ�bH�L�Cc��Qw��fB��%�o��\��lv�:��iR�L���׸U%�Ð1�<�w�?���8�� N�B�p�����������8�7�l�^�E�o�r�]�^����eH���>r���v�G���Ȼ�tɓE$��ecw��e�ҭ�hL#k� T�V%`q.	��(s�;���11�h!G�@�k&�B�#w��vW�]e4��"�fB���;Y�ކ�m����=~$��&�ߜ��^�bp��ȸ���9"��B�����N_���;::`�P�9q\K^
�G͑͜����«r��e��7b͈ A�O7h�N�Mz���kzFħ�}�4X/2_R �˅��jA������i��r���&�u`[�*�}�҂��FX(�<�^�I�<r/�z�%uj4S�t1�}aQ>�������Kw烟ЄG7ڤ{R�9� ���0Jxk�0�*F�Vc����ƽ��{�����u��cе�x�R ��I���t_�ů��_�Mg[46)�����#�}$..�7o۽������id"6���ڒu$b9�{��7ܵ�/r�S�Kz#x$������������4/)�{��6�TH�B�n�~nܸᶷ���ݻw�}�����`�ID�Be7ݘ�_|��p�m��q���d�+���0g$�Y���5�3�4�b�HaD<XUΉ�0X�(�����gx9v"���W�dv�rY�d�=j����J�	٨/��6�$�r��˸\`�у�ܝ��V�b=��T��&�{�/����଴�VKI���ݶ���&+x��so�}x�w���4��E\ �G�)�3�Q5a��"�)Z��zY�/Q�QER+���now��Ę����6HŅ(�H�v�&_#�B�k������	� ���G21�BG^��W_}�]�z�c����]&@c��D����̌)���,�K��b,���Dp��&�g!>	��A7���@j�a7����Ѿb\������6򌩣T��խbS3�R�	�?�����|A����g�Tߔ���61� ��������L8���k^�oNbv�<$}��M����N�Ѭ*%�A+h��S�L���3/�J��Y��ͣPd��D0PF�ʹ�Y��u������N��k)y $I��(]�F�,8&����w�� R"g��.Ȫ��<ƺ�9x�A�B��7��y�i��=b��G���O�4���!��>g�=�9�1�H]�1�P�q�F&�,��j�Kz��n��'�*Fe�b�a#�����������\��ۏ���N�p�����U*�:�B�}R�u���y�#kk�EȺ��[������'����Xe"�*�Q�-6����ߑ��UMbU��S��!�Fc�����L���X�s&z�QÃ�0�ge~�8b�̨������T��ZER#j�n�p��Q(X��|���l?� O�[���p�C��6�Ӧ���*��1���DY畬�r1��W@�H#7���3�k��ȳ!��h��R���;�;�~�F,U� b�/��u�ukqSx�a�ŀ�mJ���}U^�Ѱ���m��7c�4Hs+Y;����CzbC�^�ԩ�EyQF��nP�hb,����M/���F#��h�N��p�"�F.�L��ש�)�a%ϢD1,����������~|�~u�9��E)��l�]1��Δ��̼q`�0$!���4Ĩ����tax"�a�LWĚ�5�a�d(P��K�/��+��.~��FԢ��E�bW�9=���J�ўg]n(��>A�'�������B��Ud@.E$&�땤b��3��%ݐ��u�r|כ^E��%� ~�Ĭ��&u�Ri�8����DZfY�
��Յ��k��rZ�"jb��<N ��Y��I� jک���Z�7����P�bo�<N��9-3Z�*���6 >Y��W�I��Df�%qIwI�ϗ+)|�y�4��js���:�ωk���I���r��S	�n㞉 OC| �
�zhG����\�bƆ�yǛZ��M��P�3)����@���'�J�gҳ,�gܓ�i]kH������È'������1�T(WQj����ڂ�����"��(i� ��R�F�GB,pA��fX���9I���.q�&-�ǈ1&vC%�C1�Vl�ָ.s��v��Î����y(�=K��5RN��"�ȏA����j�g�9悢֍��_ 8'��ؙ���̦����wNfO��I�4��~I�F��|�߱��l[��U�z�(��5�{#j�(�qQ��>$�8j�5y�\"bb�&cU���f�4Ć#�c�C9\ �L���룶nJ׷1�gZW4���w� ��1�r#�}��IE�rS�c+R/F��Oo<�&0x?�(+R�H�����=��s��]N��c�v�8b]V3z��*�dځ��w8�&Mhf�R��?�a�޵ٔ�@����Þ@8.�K)��lbu��.���ͮ�\�)L�IX�ˉEM��{�݆��ıX���.X!G΁p���
9|Uܞ���V
1Y�G���_ �A�A|�Eɺ^5A҉�H�.�Bm(}e�^�\�:�Hb�X�r_iqQ�{A��u�M���t�-�P�ԕ��qm�'����Z0.<F��\>����Y��G�
H��Fb�^]I#�U��\	�o��E�e	�%�;l"��2���d���gU`������jD(6=�B^-k�$���L:��`����6fA���]\�ĵ1V@��տD�02qa�H:s�C�c�j��#����Z2��C�PѠi�Ub������H>+�1N\Qo��i	)E��9܎
p��U'�LaT�}& 
@���PZ�J����ڐ�G]�
���n��"��zNQ\�H��F�Y�%l_p=��Ok����Ym���(�]�pAt<p���y�.�"�%1���Tv�W ̅�D(�z�U#�@��ȹRO�d�f+�bkE%I�)���*6.�{����� ���H�f���!��X�N�q ��#>G��/�9�7�������GO�c��HD8��>m
w�֮A4�D"FmI2x�9k~튫�/�ĲU
��@�����?��Zq���ř�sL�&���5߶k̗?�m��y��_���o���P��.���b���(�r�W_�]�t�		�O�M�㦖����_�%w��Un�%~��������y2v��_cn��36�P���Z f��OZ����p�/_�5�nx~���q�nllʘirI�n���(U�0n��Kݗ������K������c�)~�J#A���Ġ�i�n�5W��j�䆮��������J��&>g�g�Y��J;j�Hל��]ߖ��e�>����}XQ0��xx�>p��l�	ӻ������{W�^uW�\��Y��0�e,�� �C��<H�����Z����%"<�`1T�㐾�A��J~�@�Y�eBl�r�`Oi�A���n��迶2,�%���!�q����1��&�3q�r+��x� �Ͷϝ�5�0cH],=�T�5Я�;wPC�z���o�
�h�0p&���g����q}��nJ�H��ZĚ)��z��'z�.�鄍Ɠ�|��V��A���Q ��E4�Hf/V�S�A��1��2����b���cU���韂$R7�<vX��:���d�|
]��(%�Z��7UhK�.9��~�tb\5�[6��[W�˒�?���`97�V�·.������p Z�IB�Y&;��
R*Dl3s�ĦK���ȁ  .,K ��"��b���sb�繩fgK|ta��C�G�B��7E��xH�'��DX�4�3#����B�[oز,��Q�!�n��|s� ��Yqlk�T��A��a	qI�ʠ�h+��' T�O����2�O�&s��>�&��鸶s��H8T��;��{C7\faF`��E\1��͌[<xu�H� �k��%�6a���'u���AeЏ@˒Q��y։1�c.�!�͉ � b}�v�]�W z��$�}�&K��Ԉ�����FV˘�5�kS�"|���Sα+9�Ƙ0	ⵓu#�<�,��Ȣ݋qo�+�Z���,4>��Zq��Hg�aQ�婚��[�����=t�̺�Hu(1:԰���H;
I���V�F� 9��2��W������J݃�Ym�G'"�l4�.�����w��++�X�Μ�-k3r�;6�!�x��U'�`L4�;�o�䳨]�mD��ֹ7�pWĝ�TV��A��gG|�5�l!E8� ����m'pu�6�|�>�Iu�%!�5�:��5wB�>ڄ9Z�UZ�9G�wi�X��δ�A�w�9w?WD�����|�	1�����o9�)�l��]�8k�\ �J� ��x�^pZj�C��C�q�E. Wݼ���U�V?1J�^��]��o��P��9�u�_l�	T
� 7V�\�ˠmݫ��v�6o�vJ�Q�NR��xAĲ��܈z���p����bft]����9�)��8�I���2�� �.�0�s-W%w:g�)�A���Gf D_+���n1�H�A��X}�e�E�J��lpF.�D���c.ͺ(��_Ծm�uq����Gc�9G�`n��.z��WsF��V��W5�Y1s�]{%L�(�v^̉쵬���dy��` �<��!ħ��p�����T^���;�o��9�p�>$�&��J��伂��i�Т5R018Ir��q�����F��i�{������'�&��TW�����|�r2\\��i��ba����e(�:%v��*�H-�8��,���6ٽ�Sv��MnK��ܖˑ4�02C9׫-/6J�����;��|�礛5���暺.a��>�]-@�|��YpwV�MPK��
�-�Э4y�����^rɠX�P�C�{�bB}WKr��za�XV��(9*�TM�Z����e�2#(�f�:�2+V�ui��5At@|�:��.��#���3MR�I[���t2�D�.(��R��;����R1�:��r�� t|�ԆУ#Y����D���NZ�q�~�Dx�1��`B��[c�Yw�=̐�۱ѣ�Kx���N�����S��	j�KdCEz�	���c�ܑyh@N�p$���0�^)�2ś����o�c��
�xwx�o��8���H&�-���h��:j��,�ei��U%TKϺV5$�]8�����"�qj7�t�Bβ�u�%xc�:*s�����e��v�$H#�rʆ��4=)�*��k#i��^O�I�x5Hp湓�BkT�F|�Se<���<�z�<S���k�]�����vx�y�jvO��%���C�!jY_�½�#t���#C3���=I�t�ʶc�lN�Kl�J�{<-+Vx4q���(��I-�,Krol�XW���i<IB��r�����xV�Ƀ&pIvg�9ͺ�I�%�%+�lK5��뭔U��\���$���S�v���fLi�Y��"�r(�����Vc،��֒��DF�\#�de�U}hR�c��![grdQ�π�M��X<�j��U�Q��,ė�����8G��%	�84�߉s"��9�^��</'��r�/l{��oP|���F'9!��o�j��X���s
R���1��։cH�ޑ�QsP�a�ԉn%Q_q���͉�r�}�B3�Z�ZT!�j���#>8�s���ԧ�v��#���t���c�чw��oLgn:�����PR3N����m����|�m�;�*�|݊fA��X��w�w�c��ooθW�(�w�'����������p9ݏF�F[������]�s��������$F)> ���h��8�l��^��{����d���U�EU���ƽ������?t��z �wH&*U�p�D>u/����t��]j�j-�`>H��h�v�{���6)oĎ'5��u�qpa�.�
��b��@�� ���"nUj8m�Ny~���'sfx:(�eU*Jz^<~��=x�1'��}N@λL5#՚ �i3=�����i|<f����o�/]8o�ֿԺr�"���K���w����sLo�X�zX�#Ttě�o��ɴ�	�Z���[�6�������/���B?b�]�������t��Mn��|�&/�3
a�-�[��Y�����������4g\k2waz�K�q���y��qY\��U%	�<��ގ���{��;ܠ�,���� ȼ�Xz�`�ELЗ�c�H�<�]�v�_�6ϵXN�)��U��WgM|���0��t�F&ĝ�t��;�9r7�%E��X_iX�b���Ieh�b�"�ȝ���$���?vSd��Eg֢󾍏�r�2Nt�]�\�{w?�����L�,W��r
�A+�\(������RO�x�!i�?qU�v�1�v����q�Wld,�����d���5���2Ă���X�M˜U*�{%����]2�8;��EB0�s��.��֔��u�	���"){;;n~��Ih�R�p ��I�dED��0�J�1��FO!�c��qJ�G�s�8�Ά��{��g�QN��l<i����ܗ�\�4잠D(0
�"#�w�̯����yQP�"j�������z�9�A4*�K4���ZX<^\ĜK����ſ,�Hvz��=�ySȿ�FE�2`a�:�Ug��[�%Q
�%�~�:�U�b���w��J�[n� �=`5��H2��g.�we�:�Ċ��
��p�>�aU�L�vj��^`	�TU�h+�Q���X ��|��.�r̜C}br���|N�/j�3��j!FN]\H�3p3.oR;u��P�]��J@X���!�Gsw4�g��r�$EjDY^+L�	1O
q3h��uԤh�؂4�@D����I!�FpI��ZQ=*f\M)���-Ѡo�6��p��b 'R ��:����驒�D���&����ld�
�0b� �1�;W���Gm!�L�� y暤e\�R���m/~�\7t�Z�zL*����`��@� w`]R@>y��3�|8�3�M7�L*�%��e���uI+8lА�w,v?��� }j1?t5�|x@ 2%�xQ�4JM�aUL���C_o����F'���#��tz�)n��Y��/$�?~���<z�R�D<tT����H���ر�bϗW��&'�!BɎ�q�j����$��Λ0d6�9�jbΑ�F��.�9�쵀��Zԭ�_��u�7�;��q,�
�qJu-�߀D�@�(��$�ٕ�yA��q���	rUA�΢�9!D_$�8`;�K�Q*V[��Zx<z�["c!�h$(&Eyi���J"!&ڰ#/UOMi�P\���/�$�Έ��{�iK�?�Zӓ�#}�Ƚ��w��G��A���t�.]��n�����*��͌�]H�	�O�8�D.�'��;��$_D66#2�4H�bK����_d!w������[�Cg���n�\��Z�W 	Q��J;D51�wU�y�N���T�wpp�sft���T�\Mu=dm@���;�*�K� �B'I'ס�Ȍ_��flmM�ܲV}2J��g��OPZ��$P!��w }��'9N���"�N߯�'ֲ8���Z���-P����4�����~�Y.�m�����~
�"�/R�}�GdIn��މ���Aۨ	��mNp�=mIrWR7K7-/4��=�pf�ݑƵ^�%D�uD1��Raٲ�BR�(i&�J��pl�I�83��:�^�9�81�@^��r>�H���&:�ظQ\Yj���tuT�DL�vWH�S�J=��R�a�ьw*��
�=Y�:uOY����9�q�B| �Z�W}Fzt�LCNHW<�#q�KK����t��Œ��o~q��h` Pâ�P�6/�!�b�VZ\_o���部�^�d��H�
y��<#)�S5+�c�IV8;'d��Я(�1Dz�y���y>��ܢ\0�ۜ�Y.�G �����xNA����L�� ���p�@6?�1��A��f��f.:!�߰/��B�Gm�P.�$N5$�.�,)�g��<z�r�g��j1��
�d�<�S%�$���D"A�'��e��.�8<���!�,4��RM��p3�hQyа��%+�X�?�;�w���j�.Nw����}!J��4�Őz���#Ql�"�Յ���꒳�h�D�0�(�i�;qt$��4��P�$
=x 48���b�cN:J\��ֲn#m�G	�d0���x�ሇ�ǆ�cX�m�[	��qG8�ߑ7��Ȓp].��>�}�ɳ��ܘN*��p]�ó">=���)� w�JA��jq��7cX=,:�doy׆������.�n�M�ݢ�fd
���3�,W���6
~)��%Mrqsڍ'x��3�@+����mďd6۔��	����p)9^`M©�K�t��y��җ�H�Jh-<���-w��5��}��E7����뺗�c�S���t�O����9
�-8�tŹ �q.��$���u�w஥tV
��3��h��9wp���L lk�s�Y�,:)a�����0kP���>uY�u\����sʄT�Cqȳ�LJ��[<�N$�|��[��|��A���N�z4�Blԋa�y���%�A�]$���ҭ�,j;QQ��
��z�os� ���Q0RI
�X�y^�\�\[��Y���P����ʃ��K��U��K/Jyu�J�>�U�޹Z� �+W���s�m�T^��j�i��q���kn�ſ��LK�5�q-!
�!�
������Q�z�9�ԯ���n����5%�Ə�Q̝a͓1�H�g��n���!�
gsDK���ԙc�P��]��"[�������R�	y�uw,�K+ ��V����SUĭ�� T\;q��i|y�P���ϳ>.��N?2�<�|��R0Ԓ]/���"�"��/�������������;��3I�V���/|g(q~����Eb5�/(��B���Xr�����R�T����͂�7C�ir6�������x��wk�j���;l�T�V����^גϏRB W�EG?�˜�%���<˓Cd2W�����ؕ\�_��n F��z��A������� �Ђ�����������`�\�)�����8���t������a��P�zX������-ū!�#ѐ��7���ε�2��p|��-,i���VL�L��}r���D`
T�6��k�*���D/��|"i�R��Ɣw�
{�-�9A��8�eDY�Ⲫ$[/�"�}�?X��F-����x�w͌P��P��y�d�s�1��q'��B��Ό7<\��n�9�$wd��⒕�e]MaH����]����кmFf5/��aNO�X�|w�Eږ����\h����(�MƆ���%�{����3�1�D��{���@���&W�ą��´_�{��^F%V���mi��F�JR�U��HN�1�g8N�E�gZ�x��f�&��	�:ײ�q���.�l2ϵL
V�{��(����g�`�ÎJ���E±x �*=��P�Lb�t�BZ�r�dpm{b�;��,��|�-�rf]'ڽ�{�JiM�"�%��C�0~��k�*x��<������`Tp�?��&1���a��,�����^���S�G�ϖ��8>8��dn����	�#jY��)�S�]^V)��[|CSta%�F�K-�о���\G��c�H9!�:I���졺h�M�2y. -(��k`���6��8�6�� ���W���cL�|U�Z�	.��`ɟ$
�kK,ĺ�� ��77t�%V}R�5���`C#���6'uA��eE��t��(5�(J`?��d� �[�Nu��·�(��4@�5���u��Z��D !�E��Z��#�MrjP�Sq>��Y�7�õ=C�k�!1R�
\ș��V\1i�;T�^6h��Z%x �%	y��P�FưxMRd�uJ/��~�?&p�ڤ�7�{u�Y���$�5��Q�ù���bw�&s&��sVܜ�-��K
��p��~�9�%�Yn���F��O�B��j��L3�d�F�W��(��i7?���ԝT�n�~~�w:�#�����[�������P1c��*Y"�SE�=�p#�[Vq ��]���poC��>���71	R@�f%�MxW.�G��ٽ�=C���7q�ͻ!����f:�~q����`/��L����#�p&�D���ja�n�$���mN����߀pf,��d�W,ciR�j�k��rN]\"ޙ��!��Bɒ��Z���I�Y[�=:BK^��u�|џ���Ɋ��Įo�>BM�{�LQV���ÕK��L6�����҉�Z�jՔl��9J�P5�Q�гI��0����V�i�����>d���{+���z�_N->N�IA����( i�g,�5��{�>�qOy-�;z暍rAAa睳�6|�tT��}���v�i7_���	e;:`�v�D�z��`���|�H��e��#\���6:[<_b8C�L���I�p�����T`cr�P��]�X"�X����1j ��3��<���qR�"f���&���p���g��@9�ح��?\=�,$��5#(!��O2��*��7j�����x�%�)�M�`����蠇"J��Z��ib%>����H�k�ьv�ç�P]�Z��`��Tn5���1�+f
g3X��xa�j�йøp�]K�|3�X�ln�"3��*w���$��!*�}yY2��e&9�qe�a�֢j��sc"0���n��,�dq�H�񌣫;b�6�E�nW�
��e�K���$�K*!�E|�$�B'%���	�!#�(� ��~Œ�%�e�5�A��=��9�2G�prb9:$MG�$��g��U[��3��p�Uj��ь���E�s�x\^$�,1�b��,�R�q�/Q���ʡo%����E��'c��)���u2��7]��nTK�BW�/�h�������ڽ���r�H���<"��gUA��gYJ�9,X�d
z0@��Q��\p*�@�*���Ð,��)^�h���z���ܾ��4z��O-�M���0?��p�ʩă9G���=D3�E@V0�`M#w�,Hdk9ȸE��Q���r��5��i��+�*�������
 Evx��M��p=���#rZ")P�ΒT�2.�y�ON�ܻ���|P�c��=���%�V)N&��hړ��Ͳҩ�d@���~\�uw��=n���x���hb�}9��G⍴@�� �����ZN&��_r���y�-�ӫ���K�w#���~��ݿq��yj�
��w��"5��P�����+�~����+\����"����� �����w�y��q�(�(�Z�D�{������N'�o��?vo}�+"v�S�bA�F|R�
�w��ΎCmjĜA�������l��0�nݺ��z�-������D���MR�|k�6����]��u�v��f��������k�$D?��&��@n�{s�`"��^W�3�o���p���j�	/ Fd^�h�i9w�������:�'�e�?�H���{�捗������~�~����w��(�[������:c�n^�ޖŰJ	@�p>?X���EiI���Dl;D�lƱ�N\hM�7���K�\�RY I١Ƃ�f�EqM ����>w�|���!r_aߨ͂6R|p�}x�cw�Ƌv����d��8��_fN�p{����6K��<�q���;K�#��>x�]�����y,BGc����ڥ��oI���\��5+I�B%�m����D��X�!E�Ro��r!9#���7�R��{4A�n�@Ƞ�p�$FAk����Y��]�*f�����I��d[��)�	%+֭�<��.�j����r����sn��o�5��O��;jc�[knmn�C�Mӕ$�ZP��D�Z�ل[�~���=�"\�{�%���c<"v��Iv�4/N�05Ё�NѲi���}x��������$�����{��u"ĥ��W~�]�~��;(!*J[s-�� [�*n�%�ݽ���Ã}"�'�c��Ľ>��G��8m�,jJ��`��	��%#퐸2�k�4a=x��,)�V/@W n�mħ92@�H#hI4��	��-rIʂ�;A\zj3$�{�S��S_J�t�QLS�[��8��N`RN���
Q�)Պ�rT��o�G����f���/^t��Dt'��(��"���΢R1"�+,����.q�w�����m��^�z�-h�٪���(��9E�����9oW�������Kߢ���7�n�����B���+׸+Q�F*�.��Ϫ���Eo�"�����I���}��I̾�"��A�`"Px矡����BQ�i�n9:gl	�e,�$��4m��r^4'�a�ꨒ<&�eQ@�!�,����b�UgJ|[[.�阮��=�tjÕ���wV���HQ/��{����}�[�r�G��n�kׯssggG0l��>����(E-~��kȊ�KYL�(����ͣEb��-�ė��U2N�0�b�����?�� ���Whg����5F�@����O��;����<_��ٹ�s�"�z�Z��Е��&q�k׮7�A��2�[F��W_��<��`��J�|h|�맺�2�&uk��J���9m�<h����DW���.����,h�;�����9S��i �೦q0X�.�+��b@����*�hE��������p��H���~��v���Hw���A�g�I�!��K~m������+r},�ڜ�*��C�3�G@J��@Vn�AL�����	aB���!�Ĺ����x<���H��v_��o����(�X�-�-�7���a�H�:ܹ��%��\��	�z����Rԏ�ƂT�B~G΁�vZ��I�T&Z׏u����S4�T�.G;2��+�:V���B��"ey��A��oE?�of�#<)pk�;N��ۙ�g0" &�������|��۷9֜5�i�<N��&ͽ��NϠ�EE���Y�\�u.�ϐC� 
3H A ��A�h��-�������GG�/��O?8:��}�pX��%�%YW%�gJ$H�$�PsU��߷��ggVPT�.�7"QU�y���^�֢g^r;�I^FK���R��*i���L/ �+�ɠի��T���n_s[ц�@��c)&�� �&��p~lD `I�D�F�(�����	M]�F����opCĔ׃!��C<��r�$�4X��5r�����n�[�Ꞁ�Uu��Q��P��;惭ӈN�`��,���7�DH|}�Q/N!9���*k��ܴ�xR�j���ò�/]Q�$�$���ׅ"�"t����N\,�3Ф(����,4�"�c��H�pŪ���5��T<ԅ�*���BAp��y	�Iī+=�D��/E�J���9�[2��I�v���Ggm�Ă*TxV��=��OV�� !�E� ����J�&�O������F-S'i0ڄ8EJ��Ԉq1�{�J�C|����?1	lDSJ���^!�Bl����v���_��$0����"�M��^�܆��
�	����+���cmZ�(�P 8��>�0CN�"ܠN$M87�������U�D�I�Cn��*S#� �F�7���ONK-@"������D���&V��_� h��,�;gC[1��ð���q.��!-pM\U��Ʊ��������)K�S��Ce�F�(�l ��.�@�7%	�k�g]�L:�eum����mj� �;�i*��p>(���%�+���k=>,u"φ���Rن�,���S��wg�<o(�ܝ�y���;����{���C��Io<����E�)'���=�2�V����~��o{"��2��B�G����l���EH�I��5����������oC���yt���Db�2�@<P&�Ɲ�6H�2,\�}��k����W)z�EoݾC�<�\#k^O�r�8���ӡQ%@]V���Vyް�H�rA>31�^EX�4��W�㍵VS�Eb�"OZj�XY�����zph�$I.mБ3�sͶ\ ZO�����T+�W�q%@�&�k��]�OW�U,
�`�s������?���x�[���Xk��Cp\K`8',]8bQ�bϞ=Bd���J���C��'N�o|����	�t�*	'���s��	�{�ؓ��*P!�T��.��>������ݹ=�+[�	���Β{���8y�bJ�e�M��g��qܩS�\��!�fx��UXT�M{��t�czޏ U}W7�+�P�^o��Y��d�%�4�Ԍ5�Vñ���]g!�[�K'7�9�3m40�U2)�ƚ=�^�iq�9_ξ�h�]5�S!2�!1;�
JC�q)�J�����������{��Y���	)��.�������)�N�+�=t���%.Q��9&9hO���9XZ6S�Οbn��C���Io6��[��FT0�_��ݙ3g��s�&���,u�{� b�!ϵQa�̸B"�a�ih�����{v�f�(!���p|"�S���.L�a�LoK�s^r`N�c��TڽREQ�6�YmP�j߭p�BuoE�4rE$)�0�Bc N����-�7�{���B*4x㛺cX���,�F'����Hu�=�w/=�"��b����db�Z*K�5B���8r�/���~7��+��/�dt����_�I�J=b�X@8�	Y\��2�{j��<[��?��Bط�@ �R/��cZɫvZܚH�������\M&�����$qV��60d�$��ɤ�'�q���ELP}���O���B�c���$ƞ�4MY
n1񴘧�V5 ��s5 y|	��>;H���d��SI5Z�]qi�Ub�P�B���j���"�d�dѼ�RClfp8�5���|�Bd��\�F�5Y����`e� ��\���DP���e04��ڏ��/��"�D`��sM<�����F >r�|J��-M<��R�.�Т�N�t��Q*��\��;�"���/[^[�6d��p�4R9D
�g���.4�7u�W��vI������*��R �^�����R�M�<�9�����9���"S�$e�r�8�JG <�&�ʭ�L�қ�<�}NT�4t�ma�P�G��}�.��M�q��X[w&��v�j]�A}�ö��A�JZ�6̗�+��6�R�Ы#F�GZKF�8�w>
��FǦ����iZw(�K�Y�
�/̾��qe
 y��S%Aobl��IKݼ�6L�Df���@����X�1�_�P��l��� @�R�M�o4���Ŏ	/vp�K�:A������� ��Zn�NU�uW�s��]��q٫�.8�B �A�)W�tIp~��`�َ�,��UP1b"�<k\O`J
�ן��R<��R[��n�u�8w���&���$�?�*7D�RI%�I�2No]�\h��MHH��bw�mal��.���ҬfϚ|m���R�;�i��e�H�a�Y<(��웑��VU��w�>��#*���D�?�f�Qw���J�^����X7H�Y��>�P
�m��{Yg��{҈H�zf��%eµ$v�4��e�ӱ�؋9rR�З5��ٸ�*�5�{��,�֊$�sc�5�S�S?׮���d�� @�8I{'�|��F�۷���+1P�#�P�-�'$Y�C�'SY���k��@�	(�� -ayZ�������� ��M���V�*X	5*%@A���N��;�3�I��2,HBa�xǉC)��i�JpN�LC�H�^V�+�:M$8��Қ:t�5�K�_n�Œh�����i
k�%&g͓�Y��MB�ăs���T�I
3FT�)ゟ�.�O����E�mw:���l���g�9q��!��%��
�:�� �P�J��.�Qf:Se�r5W3KϹ(�PVp�%R3J
��t�x��X>��i� S C��rR�D��DT*um,��ф�sj9�|W��Ҙ(�\I5�s[�";��&Ϯb��M��}2�'��6�!z_�' �o4&/�d��]�-f��:Ǽr����y��y�$Iv�YڥZ�|�t�^�n��礱Xe��<+�]Y,Q��>�� �ָ���A1U�w���;	ۉ�	tVC�L	�Z�l*1aӆ�m':[}�����D
��z|ZYȷO�.�jI�u?�抰��Uj��U��^�<��`��푔���4
�D�)7��Ia5 ~��*��W}"ڕ��`S���oT���vE	$�)���v�n�>@'=����Y�������p�,0H��|[���R�c!XxZ�L�3�(�o�x�
'-K%��^	-iU���Hˬ'�"�	��{���\]�fa�A������V�c*aX+ A�4n
���&�L����ĸm�TBzuA)ʘ�Q&�n�Ƙ����:��@B���f��j�%��l�Z��BO�Gw�hmb�5�V[b�˼  ���_����|��d�bJw�≶�D{h��D�k�f�Al��iXoڐ�p!�	��P��@�R���	���ګ�t ӻ߯��b�\�Y�n*�WL�l6Q)5s�Y�����I�@�r�է����t"'S�ED�Ot�F���;#��4�/��V[PN�j7���Rg��u�
%d^Z;�B+ T�d\�BE��Ck0Wڜ�1$���-�G����T�{F{�y�/�6P2YK�1`D_�ז�Ʀz����
�ū-�Wt��U��Obuy�-�͉�q��Z�ۈ���Kg#4��*�U�E"���w��$�Ύ5.&���
@��*w7�g�9�F2�|�J�j�+b�X�#�v���0ـc�qd�*��,/�����R���@J��= N�?���g�J]���e��>|��w��M.0 �7��ᾭ�����رc�!n̎HiM�eY[ˠ���Ub���f������"oka�羶t��͓��^��1���b�O�b�m!a|�ć�/MoY�v� 4�*(R'�:���nݺ�]�L(�T��婕?��녰{Eح��l��#�sV*����z����i�W�����?~��޾������\��tZ][#������oNTw��,d�5��ƻy��{�w܊�\N�Þfv���-O��nbr��Ɨ�"e��mFkr���M�����{��ܛo��|I�~Z�p�����~�p�;�~�7�A�z)��P�NHh7Ӎk7�N:�7?��HG���a���$�~�<���7��xf 0^ d^�������$���GL-���0]�������W��!�����
��D�iR�<qG�$�t�,��Ek��%�*Qenm�Պ9��8w�����5޶�<�e�5�I����g��{.�߭(�濢��� p�7�_s�?���Q��%W,��j���Eϝf��PrzS��&�H-% ���iqi�y��n��2O�g�"~7b�#Ԓ�z��(�(.5�$�0�=�zFp�o@��u�5O�b�f���A�nE]�,���o�ۙ ���kc���s�y�W6�-�u�@|���4�qaN]]-�HbPE(NC3����c����Չ(��t�$���~:qO���'$w*4��as�;�ҥK���u�qmĎ 8�:�AF� �KCwKs)H=YP�Swu������Uԃ�Db�n������S
z�`y��W��)�Ɛ۸�I�n
��sgVÎ	�aRš.�����f!�i����7@sJ*O�����	\��T�`�ᾄۊ>�6e}�n0~�����U���}�j�xP�Q2��o��Ћ��"k��;._ lGv�@����J/!ۡ�֠ǾL�Ӓ�P'��y�*��-����z���<!�&@�2�<��hCqmrj�0"l"o�C��js���L�St׬�P1/�Ҋ'��)nZ�삔D%k�}1Ŋ�,� �(IZ���\ <}�z,TX�I�âF���h�o�U>o�hH��I��'z�x�f�w��3�;�h�K� �p�AÝ�!m�qDh����I���ج�u�	p��� � {/��������a�D6��-���<P���T���Z���"~��I7�w�����c�O���2�~�����h�����@�N`�?�?�Q����Ϊ���	����L�n�ƥ�\��C�G��\�e�dáU���b	�0C�����k�����e�.g�Jf|��J�(n�Et|�k+qu�e��;�; �j�A�-�j�sR$a+��ei���	W�_��m'>N��/�k�1JH�K$s��	Z�[Jb�%]����괬$�Lb�֯�Zq�s2}f��V̪�5��Nv1��z',�Ȟn��"�V���{��1�L��s��$��3��"a��J�(�� M&�j=k`���u���r�-�/8��ƞ&ݞ�)�9�E"�e���M��>_i�7q'���+ij�3�a���Ăѥm$DWK��p 	4K�ɼ�����E�ܭ���-?�_��K���(�� ��j
�jh)1p
�����!^�6��Fx5��/���);�[ZXvs�g��{Cr�J�'C}�1�� � ���BU����P�d�տk�x�c�A�;mm7 �dy\M�D�q�Y��[,h��-�=���ޡK���["�g7�R�w$�r:.Ku���`�k�ڸ%�F]�:�Z�t�K�zͩ�'��b��\(���i.�;B|~�8Z*�ɪp���x�2]��RCQ���ؿTQW	��U�e��f>�g�H+����/P�Q�h|r�M����B�	vu��
eˊJ�I�'B�I;�ݵ��ʹ���HX�b���Ğv RX8�D_Y�@�v ��ǋ�<�1|����{k=��1�K�$D��S��J�4"B�>b,X�ӈ�V��\��+�C�PS���Q��`Ҏ���zl�1=A;ͣ�@UT;���'cB0�Z/�Z!đi��e!Lfj=k�U��a�O*��d�H�
�8,X;ƌW)j#����I~��6���i���C)�R�\�f@��k7�L���`MC�V�q�&���E.��a�2�w�Y�����:e�Vjh%F�O��"ӞU�CR{Z�Q�E���4�
ϠI��n�0 @�bG�ũ"H�n��.`���$����W10�PSԮ,��(�mw2WY�9_bQ�l_{�u��,�b��:D*ͧ��A��(��b;C��{�tc�~��z��X	�R����%��u��NW˻2ơ�u�:�����4������fI���ADؘ���D���~g/����B�LQ�'�VX�v�i��$�.9e!���PW V�:T��a��(��H��1�F sm�������8_G+Mu{�	�W֭I�}V�3c��0���������(3���\)ƙ���RUYzi�#�Gr����`�Q2�����g�+�G�����Z�&��z� :���K�˞�O�f��yΥ�Q��xSx�xS5Ӥ�|ȝ{���	�����a�m�tN�{��Q�qV�b�G%�u�ZYD�.�<r�4�MI��*�E�<�4���;��¶�}�eژmGp%�!O?�y79�j!�V0ବ΁�S8��8$O"	�E_)Z[���O��/�z���p�!�VC�قeы��y�*�� q9w����ԟ�!fd�lkR�Ӳ�%z���LqH�(ϝk��D�筽"*��Ô�7i�vQu ��T�D}4���1����IH���������:��~:p�U��M*�{��R���4#("��f��D��AˉG�2o�F/�-�!F�z���4yi)����敌�Ė��y���_���Y�� �C=9�D��"�8��I�}�X9#�A��Q\�%|��{���&uJn�,���..E"Y���qݞ�>`���`J��Ǧ��I�'�,��p%�!$��s�v�4��6	���?�T��%h�j�"�%�o���*�l�H8B��?��}Bl���f}�TEpi��ß.q�\�Ka#!���`e)t���$�����!�/9:���y��76����8�b�3�φ0�С�LUCם�S�ڕU���"���f^�^\e�o���^i>�z�A� �oH�Ɣ|E ������L
��-��F8���Z�m�mk��ܘ&�Y)�21?]�&r��LE�ğ�H$m���D,�N��w2qg���4ؕpTM�A�4�[5����r��î�$tY(�z�&҉"o�+l�MJ��	V�t<Cw�v���w��� ��Xmj�l���3�N �0l"E��j��\E.z^�]RjqM	���X7�K�{$�R{�����ڂ O5l���N x3U:I*b���$1[�D2�h|�Zѐ�Jtq@K|�\v��K��#F��%)FBH8\�����tKE�PAU����a�)�R5K�vU+2��p��i�^wj��مaQI�����Y5Uo��za���u}0�����F�D\��4J���i b	{��nt�A��s��"M��w����7C��� �Ep���bm�·��9KYm*=˞я䆜�΅�������8�պ3�
�MD�~(U8����t5,/VZ�F��e�ȷJ�Fȡ]���D]9$K�F��s�T��(<'$���8o�-V�fD�K�R�&(���3�?8\[:u������j��z� G��e�FbW�\����M�1��g%�>�,�*.�2	��)kh���C!�kJ�~?I�rg���e��
�-[�sRE�Ci�[�Ȇs*�팮?*J6.a9��BH�O��-�܆:yk��OU�Td�^'�833�V�*����^`UUP���ѻ/�̅B���	��(�1�J��a�kΪ��T�c԰zs��؏CcA'�����؇��K���V�Kr���v6˖�"=<���N�������cKu}��C{�,�Ǧ����#E ���&Š�u�n���:Z�����Fdi($	��I�̣���y�،�_�	"�ӯ�oR@Q��!Q��y��9�Ī�_c���ԔZts�S �ԓr���9��=I�A�O�&��3�t@�@�JWn1Z��\3��0u"�mQ������,TU�p�q1���:�"��-�a�[�n��Se(B_����ؒ�c�ė�Q��2�R��w�dl�t��n��6T�S�&r�=��AY s�J�>ٿ�#���R�#ʄ\K�Y���
;��%�+W`D��m��XL�/��J3�,�!��$y����M��8��j�l8E͸�(�a3IJ�j�e(Dɼ�OwS�+�P
u����B����u��r��P٪Rߠ9�i�:iȬeZڍ���l��G���,�aS��g��u��T�p�����Ȏ��DFr���n'b�����T�g3s�PlY���N��	W��~S�t8K8F�L��xɩHS�)k�L`�ε�T�& �����B����8�<C��hZ���&� #�"6��PIl�i�ZoY7c�d��W��?�i��ɞGb�ޏq;��,y��hZ�����6V���k]�̿j#߷<c)&N�C��N�M�e��N`l�.�yՁV���ًD8vXPj��)_�.`��}M*2�������d@*_�B��)*�-�,�.2�4T�K	�IߺBu��p�ܑ�J���~�J2�p,�>�*I��o��g�W��Uh��k�f�K�X��d��JY�$��Ad�2o�8`��j����2�Ӑ3��:(y��:�;MO3��HS٠��bE�۫"�J�� 1I�q8)��~�ؗ�G%��� ]�7�A�KL�]m�Y�Pz! �Dq�Q��ж4A��@xj�z�;+�U��{���V)aC�����~��>h*��e&-=�Q����_�O���\EQ��Q�,�$��W�j��>k�VW����ySN��}79��D.��zđ��IV&^�b�Zaz�FBrҁ�:O2.&�;�7�#6T��=�=�}�Ck%�,�AR������;2��ֺ�aN�Y��׉��,q�[�X���f��Ӳ�J���vV�B�pia���@��+ᵊ;�DE ���Z<�;D|inã~��C��Ƣ7��xӇ�u�o^��f*z�Re"����X)���9��I��g��j1�y3��l�O\�|�ݸv�E�)�S�5WJas�	ʊ=�Μ{��^�ܘ�[��v�!nɟ����p�ϟ��gǬ]��ΞuO?�4�-2]B���UQ..���f��r󳷙�C�'�����}�1���/*S��-\����R7��٧�Nڲ�A$��{U��L+�X��u������,���`׮]q�/}�^kPƑ�*���¬lDZ��H�w�>�*V���?xXbE:�z�M���c����+��_�[mq��5��,Q���	r�"GB\�Q�R:��=΅����7_c��L�%7�����^�;x��H��Z+kK�n�լ@��}��O^|���?����=zq8������K�@x�(��@�3�-Rd [d����k~S^'���UB���Q�X̵ʄ�T��K���-,���C�f�(��EM>��		��s�e�n;����uG �y��4��J�R���1rei����!�kIIVv��m�ҺՀ��/��n�Zt�%'���J��xu<��޺���v+�){!.	Hz�Nx���tKH(���\�R�
��f1#���ի������0��-��P�B��Ŵ�������<L1�M^nߺ���;�|,%�)
f�~�_-&�)�&G�����p+�K�ft��%�ih& ]DN�1�uʕ=� E�-.�����s^��5
�����f��.u}���P�C�E�hK����J}p�a��i�H*����Qt6��f�K��'%!���h�D'�O,�X�tZ�_}}���]������Иy̖+{�f�٥5��M\GE�X��D	�kv��nk(F��5e^�$��nu�	sJB����� vN,��80��A0��H�<���V���uIսy�,��L�ts��0�ؓV*���_�$_�Y=�R�<�1RC�}2y>���Bpsuႂ��(��Ui��6�)-�2A̩��P��`V@����e����F?Y����0M��GS�iS�C�J;9Ϛ����
��O'�$J�ۯ��,[��k}� (p�:���mD���C6A �~G+YɂV�]ZR����u�:2 *����Ї^�)׊T�.`�p$�b!�V@|�Q0h8����ie�ԍ��t��I�\o�}�cnii���B��Z�#��G����,��	��� �\],��YH�!�z���C*�JI��ķR;�鯆$,�0)�FHp����zx�D�	-�r�7\3kl��䦉ϫzy�ML����Qj�a��TFj0ȩ���>hְ =�VI"�ʾ�C'���(�� 3������pqsSKuNӇ�$��,e�2��I�h��'uWR�	�� X��{V]�A�����|���
[��D�?���e�t��d$��-�M��Ƽ~<����p{��\��fԚ�vpߴoJc?��c��.8����52Õ�L��\\F�,;	�YY6Q����kUx�.%@�K����j����A�.�A�~�s���(�`J���K��e�KӾ������J7��;+����7{}t���%��Ϩ[F�"}��e9�a:�KIu��Rs�RQ�R��&^%'X�]�c�3�!m�Kr4k^��e����?��T"��*zm���@�Й�>R4]+�`PY�	���� Ѫ��a:=Y%�ϴf�IK���%.�����i�HkX�͐�R�����Ma����$v�Z5�4X�Zaa�q�4�"�9���&ꇻ]�w��M4�� v�V��{�R��O�0��t�,����ĳ��]R,�"a*�������#��$�M��� ?]�TR?�G]��
@�=��
8S��ZrU�	�E�8*u"�� �Ŝb�����&yT&��
X��ʠ[��c�P�D*�b#�A�c�h��C'�'��P;��;��	뽎�kD�#oH�4�����##iڇqpJ�R���q���
���IH�>��9t{�[p�%� ᤢ��:��� ��dN��*%���X���B�-TܰN9(eȴ�O��9	NF�~b��|�Y+���@�V�o⧿���)��,}'�f�%� ��~��-�&Ao�z&kZ�DF�OdCkˈ��k���V�x��	a
.�a*���$��
?����־?5Jy ����ݓJ�@��� ����5e���E@��WO(Dz���
����3��#�����%�� Z����DY�!�N������
z�5�xcR�x�]e;�d.Xmܬ�RwWO�Lj���0��Sr)�D��3� ��BBO��
��N"ӂ{8�����!vP)j�,�ȯK�;��c{|J���7�]�-ѽF�Vx0'3���5��]�k�抺N�o��Qì/�S���b��F�lM�kF7R��,�fxB�k�b5W�j���9Ssa9��-#Y�e��*B��j���J�$*U��q��(5rk� �_��K�k�A�Uw[�g]Ʒ��*�FV2xL��o��_}(��Q�9���ysMb��7����VU��2��!|.8����V��g<QD�@R[l����lI
}V�����{AJ��M��9�C������v�K�$۫On6>���k��C��B�K	�5�ol���R\�I��Th�3,:rg��'幘����2P��Zf�6���5�+��Gˮ��;�cccfx�C�����,b��%��tMA����������6<��� h�k-�����%�x��6~�`ya4XZ���g�=1ɝ�������%:���.�W;]rP��yn�B���*�c���Um�b��?t�(��̄�Y�N8JƝ��������pc�>	�����	c�	w��SlV�&�K`]p�2nZJ��;#����C�K��T�Hi��kkB@�-������>��l�M���ּE{��9�����������r�4�~��jm�B�"r��ϱ�
w�|��i#�`���c�Wܣ��g��H�Hz��y��ט44�<����ˠM%d`��DP�%3�YJu�=3����C����H�<n���J��ꎇ�p�@ŷ�5B�\�f'O>�y,
A� k+4l�ԨI��_�U9��<V���&*������=��
�֎��v��}�Hd�9U�b�bٶ�I�U�T�$y�}��'7�O���10>
�/��`-G	���D�#G���`��Su�꾪��ih�*sZ?�y5���+kh�4ꈄǃ��g+�ˠ����T0�i�aUFsO�fx�8�ۈ�Ƃ����^ľS꾩��˖�Q�cu�%�G���R1 ��g�7W����Y�$�,�1b�B��cS��Ĕ­�t�\
d�����Y^Vzm�~�ߩ>5'����G�:�r����
�$fq��蝊l��Z$Ò0z>qVפ�����K��v������[[ʷ��R^�1��|�MI\��i[k���O��怆�T�wU�����vئ5�%5���A�~4P�Nm&~k>#wI�L$㭯����(9!Yf���n��f��V	�RDE֖$��i:5dKSm���`�ߚ�֥8/#N�����p�e�:��yN��«0l�b��ޜURtK�)�v�c3��FI�+�YU�;?v�>�*��t�;��J۬��9C����6o>@�$��v�?޽%Tb�n�~�{�rx���
�0�fzZ��Ke����ҹed &e$~m�$�)��=x'p��eVKy�LՎ^��>��A,&��2�g����y�iM�f{�LU���uN�f���IՄ�V�J3�j=X�,]�����qEMR��{���D�͟��H�s���"D��i������ȅ�@��!jX�[v]*��ª�SjcWDDg����kyUaI�u��<���AU�W����⁴{(��2�J��k$����I f��ؑ"��X�=xӋb�1���l7>���(R��٪��l�Z������:����D���1֬ѐ`q볫�-e��M������ݗ�n�'����*ݐ�ʨ���L�}�h� '�k�0���b�/�Q:F�����w)�I*F���S6���k��|�b��τ�mK��3X�sC�~� c)�w��5�IuLcđ�n�D�o-RxU�v�Y4�aM�\d�}�&�I��J��&�,�dz'S��F�]6�27���B��Z�@9\_ ��r��^��3A�>g��ITA�M��R����w�=�1�����A��$5(��CU�9�wD|c��v��r1��>���4�\B�õP�F�T�+#�@�:��s?��"�c�c��p�����ȑ8�]6�e�A���r<#�?�_"�٫*T��W=�z�u���T�T��	B{Ԡj�����bY
{v=�-�M��,�P�4�r����(�~=YI]�)�62�ߝ�.���-��Lf4�dZ��U�!g��K��]D�V���P8Xݕ>�z��:�}�1�;|�y����^g��h{3�i籹�i<Y��Gp֡�����VZF�έ?�&���3�ϹՑ��K��p�-����0�c�LFyԳ�߽��lf��!��<�-̬�M*���b�^UՖr7����Q�Z-�jX����E��v��E�`�0���v��n�7"���Q�5�HH2�a������<C�-�.���g�{ſ���FvO|��O��;A|ޒZa5���r�_��ET�?7�|UE���� GQ�Qܓ�&'�ry9]��2�.;;.3f?7
�ݍ��a-���q�9�r�S�M�|S~��a͔����7�k�܋�F�k��(�>s�����`jh����94щ��x7e��GY�w;�FL|�Dt?FU|q���m�sj���c�� �:��C� "y3ǎqw�϶r�Q��f�z�����Y06���K4`/Lq{_��;7�wk�u�&]���"������9q��TYܬ�1~��u�����5����s����6K<�bv����`�mb�����M���ǐ?l;w�f����Oӹ;|����׃n��"k��؆-�a:��6"���v��f�f��_�Q��Co��_�"k��r/u�5:�>��
|�Ǝ��M���bs+q��t#���k�ʰۮ��*ɿ���T���6G|�j�q����
'׊q�� J����fR[��������P�n�0���tȲ�l�u�3���<�k�Я�b��c3���bnh�꽖U��ʢm�r�c��emP�����z��|9:�'�f��F�Bp�h�i�F�E���ة�c��V7>DHT{�� �9���C���-W"��������\�����{�n�7��0�`�cs��\.��s)��jR�
w8�hC`����o�����Ԗ��ư7W���P�4�-�pV̩��m4j�1�u� ��N����zTQ����g���ؑ���ceY4�&.�w�ƨ���!C�=�ڻ��Y�Æ�g� ��a7A|�YUe�����u�����r�c>mBN��=�ݛ;��c�qO�[X��2�O���a:^�l#x�(bn�j���(�2|���Z������7��g#��	�'T���0��r�����JCZ_o3��s�X�k@'3z�mul�D*mO&i�%w��ͺL位|X�u�����e���ς:�	n��n�{j4m�1��d3���S����;�d�ٵ��&�����xr6v@���G��Q�O��ח5F-L��o�g�>>�n�ݽt�{�0�rp����yx�qwo?�[����d��,�����:v^m-�a����9����a�������UňՌQD����A��1��Qj�(�hԈ��\�8���m����
���Ɵ������D�o�ܣ����b|�Q�!�o7�K?d���or���6���[��RE����֭2�Mn8���!�G�����Ol����G-��u⅍w�FbsX���a�&��s�~F�w�{��m�I���|̨{_���݉*���z9lC�x���W&''���D��l�q�ɴ��~7��:�h��^��+���^�?��Ņ�s�ҧ6�%����7��0/����E}.ܨ1j#o���뽈�,e;���u_�������]'+4�u��:r�����������*k�jm�cE?��ws��wl�����7"�Q��6L����u��t4�����FcXǻ��h�K�FR��qӱ!���=����v���J�e��χ�M���a;N������3�<��t�=äI`6�PRv�R 1�����YO66M�>Æ��W�V d1Z%�����"۴Kw�<4HFs?� �6����������;�Fz��5�A�$t��kڮ4�O|��6X�4�a?ܪ��k�k���=�Kk*�o1�S�8�8�%M��Ȉ�mʊ��ψ�Z�#LS��u{��a�Faۓ�<���K�)�9/N�ح�^����b�ݸ�?��ރ��������Ū,�{�?��v���6�ݸF��5|c+�~�3۝� {G�b���th������ �b��1�V�Sn��155ſ�����v��}yy�Y��L[>�5�6�N�x6|��������"�>e :\�B#lKka����=�ms�6��s6�k��_u��XM���c��L:ȳ��y� �����޼iDh�k��F2�M�T6����]���ẻ��k����4����1?��;�c���7�&���o,&�_/b�H�tn���Z�l���l��ZFp�H#A�N��(�t[t�:��z��<�=���F�8g|��E�f|�n����)
ڵ�;]���}u�Y���6Zڠ�\8?"�����
KH����ǣ=9j���O����X���肰X�j��jb�n��agβ��hs*�����?���_<ןu�16e�z�q���W������5���	G=��_9�o�c2���/�l���IRwYg����x0v��wm�r�� �:p�@��f�K�.Y�N���R%E+��A�;�b�؄����O#.#,��������&>�i��=���te)-]'&�I��Ȳi�}�F�}��(�zE;�	a �'''�u�>���黶�k�z�/�u��5���"��&IЊ��wW����kmm�s
n�����%���ec������axx�?Ȝ�-���V�=������Ӵ�(�Ƅ�}~&���I/J����Y�����N��A��hPe���h���y�ꫯ�_|� �����;đ���ݼy�nbBy��7�믿�	�җ��;���쬻z�*ϳwό;{��{�7���B˃�_�[�o]ciqE��~��izz���W��=�V;h���=�Æ�|���3=�{�9���<�������~�~�_����̹�����$�k׮�wϿ�>����x=��#$Z,<�:��?�y��/<���F/^���9PW !��y뭷<wwG�QQ[E�T6xm�%N���&�t�{饟���{�:|�?~�}g�����9��˭��mw�cK~�Dz?-��n:���w��i��I6VU���@N��8�?{���~^����:czȿ�*�q�q�zL�&b2�H�=�������Rt*�p��@l�^�\w�̺7�x�=���Ȇ�0��+%��3����GN<L"直�y�&�o��x��o�k^��anX6 b��������/=�M�����*�;��7��w�n�p~���%��g��z�a^��?�w����GQ��}����_z�.'AB��<LMMs���\��N�:Ź�u�;x� �su�{�ݸq�_�!ε R/��6�E�5���я~����q>|�=���_x�K����@�e�U�&PX����6����Wl�|�'�M/.����ys��m��׿��w�q�����az
�_�*'����>���ԯڢ0/,̻��׿��qv��|��c�K<�x�	� m6F�����������]��3��5�Ϗ{ !�(��X8K�l(�Ť��b0�\n~q�MML�۷os��,�<�~���ک�����N�8N�ѥ����t�z�/�������Ƚ�^���{�x��Ӝ�"�.���v;�f)�@����}J�=���7��>>{��7��]��*ظ�h�Sq�W�^vo����ȯ�Ν;�����tٿ����
��x`��� �����Fu�׫�ꬭ���.���[�ka!���5�|aa�����~�����u ������ q��L+�]Y^�Baa1�gΜ��%��a�Ο?OB�y�5 r��������������݁C�9��#���?rO>�$u�K�0'�^x��C4 �����!*q��k>Ä'^�J�����kw�pB��[�����@_Z	������{��������w��F������ַ��^��k�H�H<'�Otф�����=���r�0�-7w;J|���ʥ�_~��/�'�Wd��]������7~�7��ӧ9�?��O8A��=É�v�*'���AGD7�eOhh�����Z��I~�{~�/yqw��-���������~��5�8�"�| �`\Dx��aqn�M���̦��o�"aaQ�끋���?u�7�4�.igc�&��$�w�y�^D�����pU��O�޺��a��[~M��=�>p^�8<gO8c�����������ʹ�94�����h4����83���Pgo����	U����8!����+γ�\q�.��߯2���%>?����zz���<�a��s��N�8������[��[��炓��Ʌ~����V�/^&Q������9��4+�3�J��<У�>�� ��	p.s��ĺo�\ &h����w��@�{=qcAh 8p�cG���8���y����q���t <Z����{��?�)��ujraXҏ?�x�l x���G�`H@�y��<!���'����ȏ�Z\\v��u�,oǺ�N���i�'>?�����~��_�H���LxpX�{ 4p$,&�� r᜝����CĂX>���Å�s\a}o��g���"@�7��^{�5�a��a��(�w�
@��hC��=��(�8E�Z��:����+��B�����O]��_��zҋ�cn�n	q/NvG����	��Y!UE���7��R\rzj�{��繁
uЃ�aca~���\���µA�����5���ԌWc���Ȟ�=r��} ��ް�C��{Bj���'�Nr!,>�������׿�E�C$�T,�?��B�H <�|�p(��j�6�ׂ�FX�%��<�_�b�+I�m��s��Inp-�����.	 ����J�����7>�q3���^x��������'��Ïxb~˽���\xl0p�\}�x����A� p�D+�&��~�=���<��������7���� ��h�p�X��\�>� ��\8�z����:<:�8�y�A3��/jj~9L��U�`ך�'=,X���qhJ�7=g��ߛ�����|p&�#�;�&[$��*9�c�=���'N�t]O`�x��Ƣ⾾����zkt�sͩ�3na���ځ,�j%�`,��ظ{��w��>�u����A ��� Fp�;�`�>�=� +�; �Vk�:�D�����]�|�=������ܻ�'ב�ܭ��|}��Eu�g�x�~%��\ԴY������˹�����=����/��H�L��XS��e,��ϰ 𛁻cQ�x�P��ۀ���	g-\��<�м���9�I����Q4v�u07Qn�����=n��� ��j��T�brl�E�_ZX��O?�$���E\zff?}�����<�'r8�9��C!����B�ȝ�7Gn�k�������b�%10�f�'�	pB��f�5�U�	�<o��l| :p�����O�%�(��3+��`aaX�ىI:q�_�}�q
knϞ�\DL�/~�����>	V��1��~�B��Nǵ���u����2<�	�D�a >Z� 6��+<�2�����e����2����c��A����3���y���=O��Ǘ�찰1�;�{��W� gZ]�;�t���nR�߾}�	�C�}��.P=���2+��:$�<�9�1b���:>o��#��?��{�r��
��]�W	��E���{�K��z�}a����z���w�>/�$,�c����H7�$	�D��`�a0h�p�~�?!.�\�D.��.	��s�D(;uM���|uK����qյ��F$Ĵ�$��` ;~�A�{�oem�`�8m�ɩqw��6��k�ۇ����p�x��O~��;;;�g������U�/�̸6�qX�àњ�\ �L����t�����;�Rb�L��h��80�I��������$�[�s#`ῃ?�&ـX@�_b�O��hOtND9`͚�����|�;:��Ϟy\ľ�����Н,�l��={�H�Pp,˂��a,���>�>�ē�~���ݜ݈ʈa�F"�Q���SO(�=1Cl㙠��{ �����-��������y��� ;Ǯ��2��7�f��L�������4\-x�5��Y\�v;8��'��1��k�I�~�������n���k_��NL��pn�ۂ�ׂ��5Y�yN���s�=����>�>3����0ݏ���qb����lWǦ��n�*�g XC���� ��}1\�ī��s�P#�l�9�߁���O_�~�́o~Ӓ�#���ź���w�����2?q���:+�t7�W^�u9O��k_���������WVū��	�k��81� �q��ښ���2��By��=�2,�m�c�a"�D:�o��Pp��]�qo��N����S4c ���Z&��g0b7�"�cn&�FXD�4�w�Ǿ������y�������:t=��f��?(-|�����`�z��o�(���؎��a�"C��0k�Fg�jgz��6>�a�	��A̾�v��s7X4�J��7^���w�x�����h6P)6]�k���z't4<ϳ�69�����c�ⵕPť3>p�a��Z$%Fw�C�Ҍ3���[tH�b|������^�h4`c�;�^x�E���*l��l6i��3��\ 6S�Al!����㻶x��W�U?�qUµ�	M �*�8ވ��~{n>"����lC�ˤ���C�&s��؈saE�l�l�Pذ�I�*ǰ�\�~R�����:e蝧��"��柙����g|���juK?1+�[DC���_����7�I�9��\�V��Fq��-"�Õ�08ɮ
���D�02�l�m�#�r�bUu:#�@<U�P�^����U�����ńi	JvO�c�	ۤ�����8��5�
�����S*�r qq6����&�����ϋ6�|��*􊵪z�2��p4��O,F����J�r�_�����ZI8~�z��
|b(�P�u�qS���p[�hX�FXX�X�4����8�����3�l��t#�8S/F�v>���t0d E1��p��sFb��4O钵V�$)/q�;��WWw����@$�#� ��u�f��ϓJr20%y&�g"7�n\Ot8�)@��4�5c*F�>0+���e��OO�yf�}���)�p,&jb�r90�ݓ$U/��A��9�ݣ=ð�Þ��m絍a�/x�g�d��:��%)F��9,�kV������v���W��;�ؾ���PKw<6R�~D.�>�cg�ʘ�`�3����̹a"�A��I VR�fM'6�ŢMN6֐���̠!1���kz��D@+t�Kw�pB�j@�˞�dt�9�ca���b}�Dn�[��#Z޴�p���:emX�9 سg�;>�ˈ�+�^���4�=i�W�����=��6���$A��r��I���\�g� �7��8�5'7 Vc抁�
aA8�a���.т�Qd�����m��Rl��E�9-b���՛[*�>j��pSۈ�=�k܏�t�qg��Į�`���ʄ_��%v��xq�^Cp:��oi�WT�9|/"�{����A�<>�΁�d� hȴ���� �?8��3�Neć�-5�h;�(����<	�Wo��T�X���Ng��g!>���=��{�f0�e%Ǘ��s8p�>���^uO%k+kM�[��O���RdY�ʧ���������D%~k� �6���D�����65F�3!�fE� J��5>F���beqi@d�:��<l��Xg�fg6P�����b��nP�AD���O�������jlw�ݯ}�k����A�I)�aDW
lG���J� a%��xl �����
F�f��� R�|��1�o���E��  �3"�/�g�d|%m��y���f�G^4����M䎪�0<��Ϭ]�E	t�7�	���kk�0�r�4��L�i5[��S�Q_�p>�A��U�̻�v���� �ٟ�E?M�n����njT2�A��B�8@t���	�c���(��� T�'0�D	"�[[^[.��x������m�j滼W�~��� f	����T�?S��v��"U�R��;���ܲj��<�w���"����=�6�n������>U����h��P�j4	����!�onp������A�[��&-��]S� b34�LN�q�Yzq a �oa4�A�?��Ȉ�k/q���11��-��>-���o�����"���|�k�Do 'U���.T���n��#�/�z�'�r[�h�;+�>Uxy�4��Z�&E-�X�yR�j7E��~���>��7o����)<6=������L��@8!������S��(gQ� G�#�HF����6��V,�aUE��8~�����9�06�y B�հֺ��]��h�cbV�oN�}:���6����k�2|a��ٔ�*a?.�XK�� 5�
�����;{�1�O�M@ o���5�O�:��o��zэKW.߹}g��}�������<�n�sv�96���I��/9Լ���s�0�mA�q'�f,���B�����4��ㆵh)�gז��"�.�)�*͒<]]Mw�����jY?�i>4J7|�`�xQR��Pq��P2��x <
t4p�n�ߙ���Ut{LMO������䅃-f�y�rg�5;{{���3�ss'._�詥�3�/_>���rȋ�	,"��<��C�@ 
ax�Z�I)(�;����6"�������r8$��&�b���<M;��χ�u��/x���_��0�c��$*߄������Ð1�J�"l��]{ff�O=y��Ν{��ӧ��*����Zy~i܋�����_����ݻ���녏��: B��:�B�|����e�w̵6�p^?�6��i����3�!3ڤziUzyR�|W�݆�E颱s/Z�K���^Ԛ��2�`8�ګ��5�`nz��ˏ�oO�x��O>y��0�E����5{���k3SS�O�|�g�����	�w<Ab]�V��)�����#������2dx�T�B�|eUfkk��G|Y�]y�'�^2ʚ��mv+ͩ�%����]2�U��Y���rx��ز'�7>��9s�����/|��V���0;?:����O�Ͽ�n:?��{���������Q�{���Y��mڔ��\G-d��|��|h���j�` s��w��vp��h�>�-7��-8�����_��N��DPy�t�ĩS�y��3/<��S["�x�9z��;���������?~䣏?~���l�0{�7��w����A������N2�~\u>�<�u���'Uη���S!�"wH|��vGq��ߣ{k��u�b}��so}�߻��n@���2���~Q�>{���:��?>���Mx6Ν;w륗^��^��7j�y{��k���K�_헓� qlR��	V�2�H��]sX	��0̢,w)��Ȏ�/6R��m�n߁�q�7l�ˆI�.>z�Ξ=���J�q��ԕǟ|�[W�^~viqq��cVm\���x,�#���a��L�w����~C����u$���*O|�	�`|jbWFzLH�;%9M;��5R14b�d~.��lQ�f�p�`X�9f�8��_ċ'}��'N�ٮg?u���O��>���_|��{��3�����w��(9)׵!����u��bo�2�܃���2h�Zf�� ��W�D�cE�^��y�w��-�,ɢ���ۡd��|P\1��jeb�/�n��H<G���减?��[n��'�[��x�_/}���<�;���H6��R�0]c�=�8���A��G�,��|��ؕ��Oj�Km�u�x L`��>�&�4�l��4�g�̪�e��ϋ��ӧN��ȑ#sn���?���o���r������Y���J�Y�n\�b{� �ü�4ߐB�N�@���>'3j�e�j����@��0pR��岦�hLGV/����bnn~���#W�N8ҟ��cfff��ѣ��sv��;�����Ct�\0;3��v�n���fi�#�%%CȻ����(�&:)k��C}��^�J	u�
����z�V�9ߚl���xۇ'�n�݆�B�p;�����n�X����j�ߩ@wi�M�����<��Z�����m��%���=ǻq��֩x�):��y#�z�J#��Ft��Dv+g�`)����� ����$�"�(WWV}�0Y?�}b��}�?n�{o�@x(B�0�/nwu�%�h���Dw��
�{%
u���wl~�]r��Z�hy�駉h����Ơ��p׃�{�v������n�GQ�����'�3�j$�#�6�An��p0��3�W&u7T�Gi6B��?�u���R���N�^��ƍ ��j� !~Q�^ZlM�����h�GHUd�ys� �+�^R��=�|:�+�*͹�Z u��,���\�Q�xo�o�>â���ⷤ���춃�U�����������~��}5����\����<�B����q�������c+z�p�8��&iX�4u!@�I/��>�� ��z]�Rߒ���okFI쀶
US�nuYZX-��������[w�y����f�x��������6����e�Gh!-���F=����:_e�3� ����f/ٝė�iU�%��L^6�c;�UXT�����V�ci���S�.]�һ}���mu4{�v�_��v }I�o�AޭB��~q�ڝ#�|�so�}a��v!��7�-�v֕0z��g�e�*�Ĳf�M_�|���}������-olK�����˿|�ҥK���ﳞ���L!�m��}�o���{X�n���WV�+i:���:c#2:�w��DO�����1O#>��Z�3����{n߸)݅�SQ���ˏ���[�����/������?p5ο����W�����9����IV����[?�Xz|�;;b�7�Z���Đ�Y�ٍķ
S�����3�eб��K�1�P.IZ��������?��<��?�{�����G�_|�s��9r��A�{(X:(��e%{M���Ÿ;�3�ό�����4��O���j�<���/34Qsn@��ӷ���?���796N��dF�$�=|�{b���^{mqff���.܏���������	�������'!n�D�?T�B�{���ɏPj`�x��5*����5�J�R�+�&��ŝ/��!Vbϸ\-��s��ۿ���!Ly��իW��g?�Y�s�oz���F9��\�q��?���~���>�~?b� pk�`�G���V�4VI6���]c�Tq���{��w��\6�y?�g\�S�#�<^�ɨ�p��cp�:��Y�_���[Z^`P�"�W^�N:��ĉ��_�:��~�aϡ����^��s�����e�s��{�>�����㫫�������|��w�?/,�=鯷�E�N 铸�%��wÆf�!wfec0����ګ��оë�p§���|Z����V���l�\�~�����-&Yl�����!�G��L///����{���3�����/�۷�ݙ�}����̥i����~������9ޙNg��/^|�W^yȟkr�a���oܸEǲ2���U� c����k�E`I	�}�>�t������'��.���:-���&���ڊ��U�r|~ֆ�硇�P�Q�����H8��������;K�hy䑅�gϭ�Z��u�Cz�m�����{��n���Nz�@x,��y���-A\�F�b��'Et6,�ì����(��U�b����Rl�~�ww'��㓨P�H��aX�It3rCϝ������X�QË�)O�G�g��ܝB���M��W�\IAp8�;�Z8�,�j�F�,LmF��I�(�����s�>!"�{�O������;�������{�sZ t0��������3�@Y�-Ęx���cǎ�($	.�c�H7r��7���-��p�5g�=X$c�	�'3�%ʠ��qC%^�KA?����`��܈q}�(�����ʴ���4���"D.^�N���h���|"���X�+��'¥b��Ik�vx�}Fؔ��+���6W�ǡ��ڽ���. y�6ccВ��v!����؋�������n�`�HTj��؈�8�{�'ǲ���V*�Px*�m�$$R!A��� "I	��+W����ʤ���Ά�67b�K�W�`8�/,j���i�ۭ����G�?ظԉ3`������cAQ��M��=�?�Ҳh-Q�j�pT*'�H�������a���·�?��=���</*P��x�w�{�G.;��i���Ӱr7���
��e��@�R��I3f������P�֣����D]�+��e���1��~Y�h� �K���QEO�K���W_}�-UQ��ȑc��w��o�F.�[��M}���?Gt�����k���G?v��ַ���Jd��a�VC��{��g�`����67FC��k�S���E��kB�m~�V�����]?I�Y�4<�X.��9&$H!&����ǎ�h�[w��Y^t/#�o�W����O��O�'�p_���	�����1�C���;"��1��+����g�Ȋ%Tź^����Q�����ҍ�-<e����i��������6G�i�sE��D�I��0�CuZ�x� ��u)�66�3�j�A�ϋ/��~���V	V_�:��o��
|��̟�ٟ����#��{��^��O/���M��I��V�;.$�y �0~ot��x�b��OV����Ԭ]���^��ZB��d������ģ5��q���k�����a?p+�[vm�A����.��X�kZ�wsFí�0�~�h�mb�0����i�e�;l�q�\ص�k/G��n���~�Q��Ӣ��tiw:O�	B(��w����e��9R�l�����x1��˚�A�:}����?�SZ����w�8=�^���^�"�kb��Y�G�E�s��D0�,���Ahǖ���1|�:����z�� ��Ƶp�q_�a�ݏ�`�g���t�~� c�ȕ� ��˪�$���|~��++�m��8������Qt�6��P[�a�D���Ė"�C�y�g ���{���5nA�[&�G;w�	���|�n  �&��,����8y�$-_s0�H�C��Df���e�B�X��CÚ��pT�{�A��~;���#��SV+(�)����4�|=���m���A��M2\��E��n޼Ξ��^�)�ҐU_�h�Rd>���������;s�4� ��*�v�z$�����=����6����1@� 2pH�p^X��B��� �<�����(8�����5@�x�87���\��@@����?8>��5# �����f����T��y�Y�^/=G�B�e��u&�@C����Y�Ÿ3w�(�H{D���r_��ЯΝ;G'��>�9rp�W��Ur38������������8-�T����b����nq^l
�RPv��2�p� '��W_�Og�z���g�C�7�7���0��
�~���+6T�ݷ�<x0�jU��Pj�O��Wb��
�
�<x��}?�D�L�Xk�V抾��*O@��u��Q�[�t�ޚ��V�]��T.E��k�O��uG�=ąa'�~A6���L�bp�J���=>��fÍ{"^����Olp⫞a�<q,���yqxۋ�c�s�U�W�"x"��+�Y�n�����$n��&����[�v��>pc��r<@�M-`�k�c�?�����99=��+��OЈq�*mh�5[����dZ�'��v�deewq>�� >��.�6���~�~ry&�]�`�~���̈���)Y�ٸ��0���^ � �z�gxp��?��1���r�E������b�02�8�S��q�[�tCp?<���ͷ^��v\̺	3�;�<}�x&��00DWz"�M6Cͬr�	��}���؊0v��j������S�B����+��z�n�]�d�V50o;k굧]�����}˴a��'�HX��>���^mՖf���X|����gB�2p�?��Dr��q�pN=z�=r�a!����;��)w���ƛ�Q�{��gh0 l�m-,���0� ��g��	#�D'��đ�xNLdbc+���8��0[Iv���۟���/gYދ��&���N�מ=�!���݊�\�5�4���}�6�8�.�C�tT�#��[�L�+b�������p<8�K/�D�
���iǸ�@#��k�nG46���������K���u�����N{>{~�7ۀ�Y��hz��v�����EJGG��<������">^�[�y�����~+�z�=LԲ���{O=�$!IX<X���|m8[�k��{^ok��P�
u��m�����BL�K
V �zfE�CB̅öaY{���7Y'��D,�(��u�?��>�_����hٸ����1W�\
ƀ5x1�!Ӥ��S�<�h����\JlR����@��C�wp�6�5��ovhL�Il
?]�#����}��'����5`�a��	'VݵkWiQBla�m[D���l� p�L8��O~�`��j�"�>d�)�J�ī-8�k-��� �_{��{���-�k>K
>����	��m>N��ͽN�����Ë�eqpv���(7��w���{2��`8��kD�gD�6nx����XM�v�����Dl�Sy0~����P�m�a�ӡ���g��C���E�^N�I�� ����+m����o�}���3mHha@dJb1�e0�q\.B�cW�C~C>�?�UN*UT��T���8eG���1B	�� 	�E�ܭ׷s��o��1��0��9ԠY���~���97?0�n]3�
砢ʞJ ��f  AY��"h*}Ybù��� ���e��8z� }o��g ��:��`f�4@��"@��t�k{\MA�m�@�9�{Bz����'~���|7�k��R��z�vdM�����?u�ȣ��	���r�r>1�ʥO�/ryO=�_| @4�� ��>߫���z �I��4�ʩh� +�G�k4�=��C��D�8>"c����A�+)x5��֩<<��W�ov������3K��߅�s@��s|��j�V�������V����+F��DFV<y�#M���Ϯ�R�O�4�F���/eYZF�����F���w�x��O���C$��i�j�È�n��}C��,h ���t9N���d��y�* 4ו+o2Lե=��c�g8&����^��4B:/z�5��r,�^�~'̼�{����������Bc��������*��"E߽A�M�~2�x�A�Ka���L��d��{�sR5�0����p-�����(;�@����b-%%�L.�:�Z��޲ӊ�@�ԣ,�����B�� z��z,�O�B/^g��=|�`��Y\&ua�v��}mņ`7��	����S�K1��0�X[�b����ʔ�UD��T.y��= O�+s�v��k�W�L��x>�hߠ�#��a9ԑ5�]�x�E���^T4��J���ȫ�*�K�Fe�����<W��F�
��J9� _�u,��Pd������?|�`�ӥqR�����xj�g�٬��#?�
��'\���4q���������`X'���U��a3h����.E܉����h�U�QJ�0�T��-�r�I�O�� >����%:3�f���8��������ېW��H�U��,��;=
��q�!l��c��#��X�ٻ��&Aof�������o�ZF{S'�|�V&�D�fC����D���0�f��=̼�*Si�&L��i�I��l�����̜X�Z���y!��n���8(����v5���� {�i?�50�o ���]��z������r˜ '��uZ�ߏ�^*k��C�O�+����l��Ç�>2�I�\�B6�C`r9P��sIv'E�����GH�|�d��Ų�&*�D�z�c��+N>R1�8�NO��l�: ��9���zs�~m�>ͥ*��������}���;bf�tɒ�� `��/z��}�Q5��Na���Z(?,�~������5��8��9��N�Tf���L!7^ߑ�{��#RQT�G*�Ʋ�	�| �(i���;� ���bT�t-�R�T0������A�7fU�~���Um[�����4�5+�����P��\��O*��b��k"L�<Or�p1_�i7ki���ߘ��j9ނ�G���6͸���7F��r t���������ŵ1�z�k�л�Iֿ���jBw��G�c���4>,�:�7P�/T�� �
�t�%K�Ig��t��T��S>L��]�$;�S�<`�+�Ic;|(�H�F�a��k�m3�M�%��<7��TM'pCN�KK�<�|�@>(� ��e�0j��ۨ~]��7&/��5�kTt�IM�
¤{c�Q��}o���y�%;�sr2+
.�J���S�Z{���x��[����M=��pDj�
��9G�М�URh%�F����+-//�Ƙ�j��v{��`D���B��d�w�-L�0����wܲ��hGp	M	���~T���*�E�(se�dF��p3�>%�Rn1j@���h�����N�'�<���f�<y.�=��h�Q�o�l���
R!`��cfW'NC�}W8<]6��T�)�(�C(]^Nt�����4�;��ɇc?��}l��u��c�s�eRj4�*�32�AC���a��Ro*��P]���A��h�5z@�ۙ�O�7T��T�����/� ��|��p}��i��o��z�y�"����HݭcX&� *�熡a~��/���y_][eme6v;�8zp�[��h�y+i��f�t�-�<>�v	tI�2��  q�[䲌�3�
���0�׶9�L�Z�걉�dr�T(��q��Q�$��aҩ�o��z!�[��B�'�s�Q�&դ���r�khOy����X"Ӣ K�%ҚH��d�	��!��ܟ��b6  �dq<�-�t���\��ڔ�H��-���q��<�_����*���p�ٞ-|��9i�X��e���I���>_��C�CO��+�X�Z�Rt)-��6���Ԍ�	�`A#O'�0���)���k?X0��X+BmO���SYɭ��=�F���W���磷`�yL�0� ~�(o����8��	!�)� ��"Of�)*r�:�P\���W�w:�
�M缰�N�l���PE2��n8BR�A	-ɭ��s��T������bӹ�2��N�"`��e�]���8�A�M�ǎ���P��x͕k���+���."z�j�iZI��HQ�����F`��.�����͜I�H�g�z��%�*���<j���I���<�����׃8�k@ � �u���С��n��?ȥ�o��/��A���Q�YMK�:�
(:.����oO��qq�����w�����ƕ��Y�k�ֆ&�s�廬�ͨ�!.�H��:ɻk~N<�أ�ر;�C���7���o<+��](�2�������m�_4�L�X��0����)߰��J������'��~0V{�f��J�Д�R�0�Ȩ�;���܂j*�+���P�Es$����K7���w��h.�"�����$哯�W�h���b����]�C7��}�㳏=.ڤ��s��^�tQ�I��9����rs�ny�5�[���������;x��x�t�T uqߛ�g���8��k\ٰ��z�f�>M�*	VY�V��\o��E��Á���$���pt����&���͌�"��4U�̀I�* ��Ɲ�^:�4b�����{D�z/�}�ŉ�犂�옿��|����,5DIt(��}����m��ffľ�{������~O�N���9���;|;�:�'�y�<���J��G"`)���ĸ@MqBעິnQ�>�дSB؟#�r�Ϸ��^C�.AaƖ H҇9v�����l�O?q�P�ϴ(R=x�݌s xbc]PZ�b������69�qϛ�PLϨFlԣ�T��R��HZ��R�h%�Q��N�Oh&���䣑����T�Nr�j|2 �е�j�E"�ǘ\.c	&!�# B�=��޵kK���뤉����>S���E�i(���!J<Y@��J]���qm���*�MRꞨ.��������j�E�O^mW�A$_�&�͏��L��
���T��@o��k����Uq���~o�SfH�E.0N"��M���Tw�M�F1�Yr� �����ϦR(�J����33K�]A4�4�>k�o��1�7��9�k�!��@_�c�A ��AO��:
4��J.��(��b��_�]���"�a"�w1�F.� �י�>ѐ��#y$��\�ڷ�Y����\�> �&+�q%�vk�1���ծ(h邔q���!=�7<�c����e_���E[UV��[=х4ݞb���;�c�Ǹh����t� >n��Hym�K�W�Eչ}8<Ќ�/¸&�JU�œ�noM�����e���҈��@,鉱S���[a{��%�4x�}�Z
Z�M>i���i�0�U���f~v���F���@=��uf�ut��u-���4-��D��	Xf�hޟU�EI��b�OMuzq:���7z�7|ʊ2;BgcB������ZpD�j@����G,][摳���QϪT� �j
e' ��j��(��Ge��z ,L�ך�M��a(I
�e]Vg�r���t�*�����Զ=�B������`�BF#]�h:h�,���Y#o�󞙞���$fR.T�d��3�[��� m^Y�1�G�G�������q��1�N�-|��:3�ngf����u~:����M�v��HHU�T5��Y����Z�Ҡ�w0+��"�}+5�1g0Н�\ �#����x��-QηN]!��)YB��sD9I�Wc��r�>i����;�@E0�R��Ӎoϴ`���4�9H�9B����K����!'�m�޶t8���u��o9�ʠ	ɷ�� C�����=�\��������̢NR�q�=�Y��&��A������J�ڗ� ��q܈�	���bN��\7pK:��ov��ݍSE�\8q�k7<�j�ͮM���5�T��$]�D��
 �8�����@���;������^��u`��#��`����.|�ї09J��wRѡ�" �:y��:]�Q�z�����rm�
D��[��e>Z8c�~��"%s9�-�{y���;L�ghf6�d��;b��s�NZL�cͫ�+;��.h���/�s��f�f^"�՝�1��u���ɳa��+K˻�;��ϋn������z�����(�c�۹�b+�X����ߴr�葵0�ٻ��oX�A6|��X��0 rH7�m(HF�US����1p~�z��bG/�8q���;�ɋ_����=���3���Cז�2"�#���O5�d���XED>8t��[;w�\��	/\��giei����s����& g�c�G�P��	j0]8WH� �Ej/����ٳ�Փ���ӛ��y��s����ON=|���#�����=hh"���]'U���-	�!
�z�؂���ێ���'��ƓO>�ӝ;�V��N	k���)FtY�8H ��/�Mɡ{a7���n%�3�ݻfE����t�QP�j����*��W��C�<E�%t�S�̱e�,�\Y�Յ�|\���p�{vn8=5u�۽�SSw�����������g����|���l��&�c!�EIJ��DɵcsC���$�n
�VY���o�/���~���ά���|���~������--��&�nt�RgF ��{a���s�^D�J)8Ȓa��R�v�u���W��O��=|���_|mf���{����p�d�<��q�`jz&��$H�Q�!J��x��k;w�Z'��	�Q�3{�����O|���O�Ĳi�#�a�S������=?77����=(�Ji��rpy��W�)���Ȁi'p���ۍ�­��ue߾}t���g6\��?�������O����:�M~[�n��ld������(NAPkO�za��v�m�{��ǿ���}��ѣ��:�|�j}�J��+�y�Ň	z}�����޽+��u����x�37ۧs�:�k�۝��i�+d�S�;���>�g�����=+����z�Tozn���g�<���K%N��Lg����+W��Nv��Y��X����?z�F�d9�Z��욝_;v���ɓ'���l����/-�:u��i��Ku�8�Xy�� "�f��
i��#�@�H�}6}[j������8����]��:��N�E�q��|�O��;�k�+�?��_����f� m��u�rW�㎥#G��M�c����n������y�嗿�y��iq���W�����˗/1J�}��<a���w?s�'>��!8Eh�tZ��w?�f]���ѓ�.��替&�~�̹y�]�A��_��+W���q�~hK҆�w�q������j�T2�-&�p<����}_y�ᇯũ�ӧ;�!��)�^7��K��ݺ��ս�fs�̚K����ǎ}�ɧ�|��W) L��=����o�R��-�e�y��ϒ���Ad�պv����������>�f��op��z����� X\B_�W+�gf��p,�	�Mg�|�bY�↯V���s���l�q-Ǳ����μ23��ÇG����׾�wLF��УԶ,y�A���߇�=��Ӓ�b��C��+</�^�	 �|���|�%n��di�S��{��H�"�n`�����̦�a��L�q�J ��y��b�
aˢ�Hs#A�{��I�l0pS�����#���IS��� �����l�c:Sa���A��cڮ�S\����v4Ѿ�	�-�4��h��ܽFZĢx���Z�4�����\��)��v;o�Zc�\-R��J���f!�c��˖_���ZS�4N%� �9L��q�GZ��2����E��� A����&��e��yNT��8��P�r�s�A��,m`��)�T��c�h������S��c4���[�ϊ�^-����F0�|(�MH����m�|�!v��]������{����c�@�s#Ij�`}QN�׫�'k6�8��6yI����� [|���i�I(fCN@��/q�A��Q��@b\�g��Vӌ�)�k�}b�@i3eˁ/M�</dY%���Tc;�q��i�pUP����H��#���������+�(�`.�P��7(�H�L� o��a�S���vvp�
�54m9dieˁ�O�{�e:5
BZB3��=6�|	���v�+ ���"��Uu�0�F�}�I�bȍ��2� 
Q� ��y�nv�٭|l��������~T����=#X��f|�qD�Ѯ��_����Q��# �:~X�{�6�#��tT�LU7xS>v��aw�n0*��dY^K�>�^�����&���r���+,�f��a�h:
�:*�J�E�Y���~��+X� ��'�kԍ��{�}�([|�'3����a�Y�]���c�
�K{(�(�/��Z�H۠� �$}��	�M���$���&
�/9o�u������m����n>%z[Z��U����l9�!p�+���\2a���\�k�+�|���*�_�$���|��x,�%�'�<�bjj�h��I���9rdl�H��DG^�e��H�W��Aq5�,&�߃l9���/n(j�N�bCۖ����J1����
�B���ٛ��Y�EL�L��߈���)���_ǉ������.�AH~YT��v�����||lz�$��->��B���d^x�n�Щ��D��#�T�e�dwk���ІzS'�) ��$	4�m@�A{ Y�(��D���5*����,�jI`�_�����4�
C�����������>h$$y�@��y��ؾ�+��r�͔�Z\�5&�嘪��\��%w!j��&�P�r����e��a�-*Uɑdl����AcEG�`0�=�W�p�>E�.3�7F[M��mv'E��T�������1�����'�=���'m߿�F������w���&L,۱y����n��bXCJ$q�:�U���k+=��
�����@G|��h���->�a <�Yg2��֧8��Y�r��>;�%Ϸs�NI��4z�j�fn��ʖ_�K[G�fxxQ�U �D�dn����H�Z��'@�W"g�2��	�->ŹV��t�-��������Q�y�4�hN��XOC��s�(*[|�v��jj/�����B�;��v�ˬ�3��;�I�a>�4v�y���j�iU�?�%��=�L ��WvsD긹��������f̔�pG��[;a@&R-xXtϮE,oG��"�%%i�������)�a��uj[�ni�������cȉ'���G1:�4�Z0@ %&T���(vz�����n����j�Y��6v߮�D���S�T�l��/��K	|���͇}ۚoRM7I�G��\KX.��f��x�7R���B�v�,�CQ��"|��_ͪ��S*[|�F���/q�����[c�/�N��4-䱱r���N��H��U��� o>�`c��N��^�� bD����N^[�$��-�~�����$�|�r- �����ouԢ?4m�oR�+dj���!�w����,N����$�h)��8�jDj]e0=*C��Ռ>�v1����״����A4��~a0�	��HB�r����S�Fl�����6R�_4�`{V�$�@�,����*riI���H�������ƫ���Z�Pץ���A(AJ���Ʊ�����H��6E��&dZҖ��]8��s=#qy�*���R��)��=/�q�	E1��$�N�L�h^�����ة���i 	E�Ֆ �\e�����"j
=�YlI�pcok�I�I9U��� �.t(��j��� &Ǳ�ly8��a]�<wA���D�':��l��21��,��k�D�0�0��r�cK�|�� ����Y��CQ����	כX�ǲ����.�"g��h�gv��	 ����:���\/A�E/Ŧ7O,�t��O-��y�Q��Zn��ya���E�ܜ^XuM- 	��m��D
7Ș[�&&T��B����^@Q�F�q%d�b�
��ډ�QQ��橃c7M:}�gK�	�->E����n��dՒ���D�42SQ�G�n]+�>zfP� ��mב���d	 �0�th&s=��ˉɏD�74�l���I��#��(���*4�#��ߤH�eҵ����]��d�6�خ��@ 7�u�|���?7�d� ��a�[4��̓"䓡�u�)��mٹm岮!�t@�x��b�\��<_���m�k�������Ońʖ_F7+�2"�)F�/˱���z�����8�di�v�]��ҧ ���<=��ݻ�7++�G�س��W�hX�Y��eˁ϶��oLOO_m6�A�|���ql������o�SS�v{�\�z�Gַ�cCz�3˽^����.,/�}lee�;?ӊ�P�r����z��[~x�С��ј�8���]�8������/������o�o�w�~r��3��q|t��?^^\_�^�zu���'߾&&T��N�<�����v�n\!C&�`=ٵ�Z�ٿ��e��Vw�Z|��v�[fW^ j}����fɖ �>4��5�ă�Ö���]���n�    IEND�B`�PK   �r�XN���       jsons/user_defined.json��mo�6ǿ���� ��D2�R�錵����!((�J�:�+�MӠ�}ԃc'e)�_92y?�x�����+�y��ο('�V�����u���8�d��7a9t�����Lޕs�s�I�l��l>:����ib&D��7Y�`&lG���(Ϣ,-�l�Թw=��'���7z�%�G�"a��B)@#�A�0ʧ!����N�:ʓUQ�z�|�D�o��/R��08����ci1Y�7f�*Igi�yG�^��;I֫�|�fK�s�	ÄC3l��yv_�'BJk��6i�mc����E�'ƾqh9 ['�J?&K���Ld,D����N��it��f��+K�r�����5n��,뼶�3��X.�{�ߟ�8�c˼j���r�O,��QQ:V���
��l6�_.���I�t� E�('�N��I�dBŇ(�8A �x�)��?�6�O��i#�9oq���G&*\nGl	�@t2����!� F�����=W5���\�ݔu�|5��+d�|�[�(�M�����%H�\B咷����`����%����:���qDJ	Do����w��Un������"�V9�@��_���7�\�Ǣ��N���F��`[܈ק�Y_�����u�a����cw�ö�1j�����)�\�x�}w��-v#3&z�wK �\մY��\�[nj�}�mߖ0�z�O8�����e��@��������/ẅ́m-�SPMA����l1wט��qP2L����Օ0H��w�޾��37�E�{����HܤEջ�E���j��pߜ�톴H����\v@Z����!�EZ�ˀ�	�EZ4�^Apg)Ң��-ԟ��S��M�1����:����&��F�\�O�n��l�mA֟ ܄��ۇۚr���%m)��k�߯A�eM[�o�/)n]Ӗ�Gt]G���5@w�	Q[ڢA8��v�-m^����-t]��.���}�ke��*�V:/���i�$Q�����$� *BN�<� �\�L#�bߗM�0��7�Cɦ�4_�_"��'�ݭ�T��ն����>o���yY���Ok���M��A�u��F@�����)�*%�>�C�TU8�@[�����BK�!T�HF �B�Q��V|�'�I	��C�ǀRi)b3��	_����՛&�2`m�YL�<[��^�c�ܺ[�WSwoӾ8�A�/�w�����״/:�P�>���v��ݙ({�o�����6C���>�1�D�Ph�JsKI	0�����2�Z����Zh�t��	��Ū�Ͽ�⢉��̓��;G�e�e�Ԗ+��CY��`�C���|R��(�~�~W����2����l�UR�aF�c-�}��ۦr}b������@{OR���mv?O�rVO�n}���d5�&
���Iq�xrD5io	;t(��7y�I��a��������oOm�+=�h����*X}��*���"���_abo!�l�'&������<��p
Atlb�*�Mtk8b�bm�hk��J����PK
   �r�X8�uȇ	  V                   cirkitFile.jsonPK
   �r�X����7  �  /             �	  images/2b66d102-ef9e-4dde-8ee7-817842500f7b.pngPK
   p�XE�U� z� /             8  images/3e05991d-8fe2-4671-87ec-9014655f7ce9.pngPK
   p�Xx[ǩ� ; /             �� images/628760d9-b837-48ba-be8e-acb7e191f55a.pngPK
   �p�X�J �i P /             � images/6a99ea4b-7804-4d0b-a50c-ccb121b20ed8.pngPK
   �r�X�&�}[  y`  /             �� images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.pngPK
   �p�XT��_�  K�  /             � images/aa07afbd-658f-44ac-9cd7-fcb1529195ab.pngPK
   �r�XN���                 3 jsons/user_defined.jsonPK      �  `   